
module dff_533 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_532 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_531 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_530 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_529 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_528 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_524 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_523 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_522 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_520 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_519 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_518 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_517 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_516 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_515 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_514 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_512 ( clk, q, d_BAR );
  input clk, d_BAR;
  output q;
  wire   d;
  assign d = d_BAR;

  DFFX1 q_reg ( .D(d), .CLK(clk), .QN(q) );
endmodule


module dff_510 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_508 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_507 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_506 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_505 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_504 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_502 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_501 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_500 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_498 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_497 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_496 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_495 ( clk, q, d );
  input clk, d;
  output q;
  wire   n2;

  DFFX1 q_reg ( .D(n2), .CLK(clk), .QN(q) );
  INVX0 U5 ( .INP(d), .ZN(n2) );
endmodule


module dff_493 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_492 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_491 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_490 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_489 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_488 ( clk, q, d );
  input clk, d;
  output q;
  wire   n1;

  DFFX2 q_reg ( .D(n1), .CLK(clk), .QN(q) );
  INVX0 U5 ( .INP(d), .ZN(n1) );
endmodule


module dff_487 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_486 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_484 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_483 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_482 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_481 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_480 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_479 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_478 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_477 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_476 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_475 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_474 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_473 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_472 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_470 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_469 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_468 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_467 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_466 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_465 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_464 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_462 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_461 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_459 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_458 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_457 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_455 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_454 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_453 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_452 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_449 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_448 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_447 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_446 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_445 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_444 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_442 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_441 ( clk, d, q_BAR );
  input clk, d;
  output q_BAR;


  DFFX1 q_reg ( .D(d), .CLK(clk), .QN(q_BAR) );
endmodule


module dff_440 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_439 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_438 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_437 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_436 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_435 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_434 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_433 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_432 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_431 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_430 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_429 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_428 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_426 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_425 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_423 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_422 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_421 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_420 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_419 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_418 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_417 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_416 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_415 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_414 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_412 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_411 ( clk, q, d );
  input clk, d;
  output q;
  wire   n2;

  DFFX1 q_reg ( .D(n2), .CLK(clk), .QN(q) );
  INVX0 U5 ( .INP(d), .ZN(n2) );
endmodule


module dff_410 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_409 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_407 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_406 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_405 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_404 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_402 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_401 ( clk, q, d );
  input clk, d;
  output q;
  wire   n2;

  DFFX1 q_reg ( .D(n2), .CLK(clk), .QN(q) );
  INVX0 U5 ( .INP(d), .ZN(n2) );
endmodule


module dff_400 ( clk, q, d );
  input clk, d;
  output q;
  wire   n1;

  DFFX1 q_reg ( .D(n1), .CLK(clk), .QN(q) );
  INVX0 U5 ( .INP(d), .ZN(n1) );
endmodule


module dff_399 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_398 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_397 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_396 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_395 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_394 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_393 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_392 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_391 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_388 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_387 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_386 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_385 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_384 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_383 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_382 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_381 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_380 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_379 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_378 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_377 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_375 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_373 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_371 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_370 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_369 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_368 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_367 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_366 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_365 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_364 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_363 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_362 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_361 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_360 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_359 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_358 ( clk, q, d );
  input clk, d;
  output q;
  wire   n1;

  DFFX1 q_reg ( .D(n1), .CLK(clk), .QN(q) );
  INVX0 U5 ( .INP(d), .ZN(n1) );
endmodule


module dff_357 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_356 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_355 ( clk, q, d );
  input clk, d;
  output q;
  wire   n1;

  DFFX1 q_reg ( .D(n1), .CLK(clk), .QN(q) );
  INVX0 U5 ( .INP(d), .ZN(n1) );
endmodule


module dff_354 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_353 ( clk, q, d );
  input clk, d;
  output q;
  wire   n1;

  DFFX2 q_reg ( .D(n1), .CLK(clk), .QN(q) );
  INVX0 U5 ( .INP(d), .ZN(n1) );
endmodule


module dff_352 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_351 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_350 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_349 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_348 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_347 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_346 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_345 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_344 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_343 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_342 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_341 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_340 ( clk, d, q_BAR );
  input clk, d;
  output q_BAR;


  DFFX1 q_reg ( .D(d), .CLK(clk), .QN(q_BAR) );
endmodule


module dff_339 ( clk, q, d );
  input clk, d;
  output q;
  wire   n2;

  DFFX1 q_reg ( .D(n2), .CLK(clk), .QN(q) );
  INVX0 U5 ( .INP(d), .ZN(n2) );
endmodule


module dff_338 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_337 ( clk, q, d );
  input clk, d;
  output q;
  wire   n1;

  DFFX1 q_reg ( .D(n1), .CLK(clk), .QN(q) );
  INVX0 U5 ( .INP(d), .ZN(n1) );
endmodule


module dff_336 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_335 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_333 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_332 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_331 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_330 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_329 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_328 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_327 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_326 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_325 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_324 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_323 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_322 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_319 ( clk, d, q_BAR );
  input clk, d;
  output q_BAR;


  DFFX1 q_reg ( .D(d), .CLK(clk), .QN(q_BAR) );
endmodule


module dff_318 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_317 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_316 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_314 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_313 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_312 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_311 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_309 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_308 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_307 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_306 ( clk, q, d_BAR );
  input clk, d_BAR;
  output q;
  wire   d, n1;
  assign d = d_BAR;

  DFFX1 q_reg ( .D(n1), .CLK(clk), .Q(q) );
  INVX0 U5 ( .INP(d), .ZN(n1) );
endmodule


module dff_305 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_304 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_303 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_301 ( clk, d, q_BAR );
  input clk, d;
  output q_BAR;


  DFFX1 q_reg ( .D(d), .CLK(clk), .QN(q_BAR) );
endmodule


module dff_300 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_299 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_297 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_296 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_295 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_292 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_290 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_289 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_288 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_287 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_286 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_285 ( clk, d, q_BAR );
  input clk, d;
  output q_BAR;


  DFFX1 q_reg ( .D(d), .CLK(clk), .QN(q_BAR) );
endmodule


module dff_284 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_283 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_282 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_281 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_280 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_279 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_278 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_276 ( clk, q, d );
  input clk, d;
  output q;
  wire   n1;

  DFFX1 q_reg ( .D(n1), .CLK(clk), .QN(q) );
  INVX0 U5 ( .INP(d), .ZN(n1) );
endmodule


module dff_275 ( clk, q, d );
  input clk, d;
  output q;
  wire   n1;

  DFFX1 q_reg ( .D(n1), .CLK(clk), .QN(q) );
  INVX0 U5 ( .INP(d), .ZN(n1) );
endmodule


module dff_274 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_273 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_272 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_271 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_270 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_269 ( clk, d, q_BAR );
  input clk, d;
  output q_BAR;


  DFFX1 q_reg ( .D(d), .CLK(clk), .QN(q_BAR) );
endmodule


module dff_268 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_267 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_266 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_265 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_264 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_263 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_261 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_259 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_258 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_257 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_255 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_254 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_253 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_251 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_250 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_249 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_248 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_246 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_245 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_244 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_242 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_241 ( clk, q, d );
  input clk, d;
  output q;


  DFFSSRX1 q_reg ( .D(1'b1), .RSTB(d), .SETB(1'b1), .CLK(clk), .Q(q) );
endmodule


module dff_240 ( clk, q, d );
  input clk, d;
  output q;
  wire   n1;

  DFFX1 q_reg ( .D(n1), .CLK(clk), .QN(q) );
  INVX0 U5 ( .INP(d), .ZN(n1) );
endmodule


module dff_239 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_238 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_237 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_235 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_234 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_233 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_232 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_231 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_230 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_228 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_227 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_226 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_225 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_224 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_223 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_222 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_221 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_220 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_219 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_218 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_217 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_216 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_215 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_213 ( clk, q, d );
  input clk, d;
  output q;
  wire   n1;

  DFFX1 q_reg ( .D(n1), .CLK(clk), .QN(q) );
  INVX0 U5 ( .INP(d), .ZN(n1) );
endmodule


module dff_212 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_210 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_209 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_208 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_207 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_206 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_205 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_204 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_203 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_202 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_201 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_200 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_199 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_198 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_197 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_196 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_195 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_192 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_191 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_190 ( clk, q, d );
  input clk, d;
  output q;
  wire   n1;

  DFFX1 q_reg ( .D(n1), .CLK(clk), .QN(q) );
  INVX0 U5 ( .INP(d), .ZN(n1) );
endmodule


module dff_189 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_188 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_187 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_185 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_184 ( clk, q, d_BAR );
  input clk, d_BAR;
  output q;
  wire   d, n1;
  assign d = d_BAR;

  DFFX1 q_reg ( .D(n1), .CLK(clk), .Q(q) );
  INVX0 U5 ( .INP(d), .ZN(n1) );
endmodule


module dff_183 ( clk, q, d );
  input clk, d;
  output q;
  wire   n1;

  DFFX1 q_reg ( .D(n1), .CLK(clk), .QN(q) );
  INVX0 U5 ( .INP(d), .ZN(n1) );
endmodule


module dff_182 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_180 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_179 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_178 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_177 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_176 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_175 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_174 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_173 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_172 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_170 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_169 ( clk, q, d );
  input clk, d;
  output q;
  wire   n1;

  DFFX1 q_reg ( .D(n1), .CLK(clk), .QN(q) );
  INVX0 U5 ( .INP(d), .ZN(n1) );
endmodule


module dff_167 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_166 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_165 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_164 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_163 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_162 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_161 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_160 ( clk, d, q_BAR );
  input clk, d;
  output q_BAR;


  DFFX1 q_reg ( .D(d), .CLK(clk), .QN(q_BAR) );
endmodule


module dff_158 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_157 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_156 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_155 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_154 ( clk, q, d );
  input clk, d;
  output q;
  wire   n1;

  DFFX1 q_reg ( .D(n1), .CLK(clk), .QN(q) );
  INVX0 U5 ( .INP(d), .ZN(n1) );
endmodule


module dff_153 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_152 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_150 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_149 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_148 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_147 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_145 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_144 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_143 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_142 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_141 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_140 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_139 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_138 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_137 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_136 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_134 ( clk, d, q_BAR );
  input clk, d;
  output q_BAR;


  DFFX1 q_reg ( .D(d), .CLK(clk), .QN(q_BAR) );
endmodule


module dff_133 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_132 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_131 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_130 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_129 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_128 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_127 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_126 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_125 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_123 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_122 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_121 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_120 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_119 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_116 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_115 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_114 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_111 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_110 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_109 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_108 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_107 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_106 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_105 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_104 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_103 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_102 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_101 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_100 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_97 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_94 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_93 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_92 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_91 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_90 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_89 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_88 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_87 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_86 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_85 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_84 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_83 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_82 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_81 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_80 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_79 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_78 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_76 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_75 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_74 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_73 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_72 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_71 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_70 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_69 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_68 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_67 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_64 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_63 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_61 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_60 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_59 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_58 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_57 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_56 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_54 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_53 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_52 ( clk, d, q_BAR );
  input clk, d;
  output q_BAR;


  DFFX1 q_reg ( .D(d), .CLK(clk), .QN(q_BAR) );
endmodule


module dff_51 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_50 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_49 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_48 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_47 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_46 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_45 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_44 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_43 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_42 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_41 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_40 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_39 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_37 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_36 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_35 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_34 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_32 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_31 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_30 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_29 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_28 ( clk, q, d );
  input clk, d;
  output q;
  wire   n1;

  DFFX1 q_reg ( .D(n1), .CLK(clk), .QN(q) );
  INVX0 U5 ( .INP(d), .ZN(n1) );
endmodule


module dff_26 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_25 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_24 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_23 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_22 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_20 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_19 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_18 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_16 ( clk, d, q_BAR );
  input clk, d;
  output q_BAR;


  DFFX1 q_reg ( .D(d), .CLK(clk), .QN(q_BAR) );
endmodule


module dff_15 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_14 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_13 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_12 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_11 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_10 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_6 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_5 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_4 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_3 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module dff_2 ( clk, q, d );
  input clk, d;
  output q;


  DFFX1 q_reg ( .D(d), .CLK(clk), .Q(q) );
endmodule


module s15850 ( CK, g100, g101, g102, g103, g10377, g10379, g104, g10455, 
        g10457, g10459, g10461, g10463, g10465, g10628, g10801, g109, g11163, 
        g11206, g11489, g1170, g1173, g1176, g1179, g1182, g1185, g1188, g1191, 
        g1194, g1197, g1200, g1203, g1696, g1700, g1712, g18, g1957, g1960, 
        g1961, g23, g2355, g2601, g2602, g2603, g2604, g2605, g2606, g2607, 
        g2608, g2609, g2610, g2611, g2612, g2648, g27, g28, g29, g2986, g30, 
        g3007, g3069, g31, g3327, g41, g4171, g4172, g4173, g4174, g4175, 
        g4176, g4177, g4178, g4179, g4180, g4181, g4191, g4192, g4193, g4194, 
        g4195, g4196, g4197, g4198, g4199, g42, g4200, g4201, g4202, g4203, 
        g4204, g4205, g4206, g4207, g4208, g4209, g4210, g4211, g4212, g4213, 
        g4214, g4215, g4216, g43, g44, g45, g46, g47, g48, g4887, g4888, g5101, 
        g5105, g5658, g5659, g5816, g6253, g6254, g6255, g6256, g6257, g6258, 
        g6259, g6260, g6261, g6262, g6263, g6264, g6265, g6266, g6267, g6268, 
        g6269, g6270, g6271, g6272, g6273, g6274, g6275, g6276, g6277, g6278, 
        g6279, g6280, g6281, g6282, g6283, g6284, g6285, g6842, g6920, g6926, 
        g6932, g6942, g6949, g6955, g741, g742, g743, g744, g750, g7744, g8061, 
        g8062, g82, g8271, g83, g8313, g8316, g8318, g8323, g8328, g8331, 
        g8335, g8340, g8347, g8349, g8352, g84, g85, g8561, g8562, g8563, 
        g8564, g8565, g8566, g86, g87, g872, g873, g877, g88, g881, g886, g889, 
        g89, g892, g895, g8976, g8977, g8978, g8979, g898, g8980, g8981, g8982, 
        g8983, g8984, g8985, g8986, g90, g901, g904, g907, g91, g910, g913, 
        g916, g919, g92, g922, g925, g93, g94, g9451, g95, g96, g99, g9961 );
  input CK, g100, g101, g102, g103, g104, g109, g1170, g1173, g1176, g1179,
         g1182, g1185, g1188, g1191, g1194, g1197, g1200, g1203, g1696, g1700,
         g1712, g18, g1960, g1961, g23, g27, g28, g29, g30, g31, g41, g42, g43,
         g44, g45, g46, g47, g48, g741, g742, g743, g744, g750, g82, g83, g84,
         g85, g86, g87, g872, g873, g877, g88, g881, g886, g889, g89, g892,
         g895, g898, g90, g901, g904, g907, g91, g910, g913, g916, g919, g92,
         g922, g925, g93, g94, g95, g96, g99;
  output g10377, g10379, g10455, g10457, g10459, g10461, g10463, g10465,
         g10628, g10801, g11163, g11206, g11489, g1957, g2355, g2601, g2602,
         g2603, g2604, g2605, g2606, g2607, g2608, g2609, g2610, g2611, g2612,
         g2648, g2986, g3007, g3069, g3327, g4171, g4172, g4173, g4174, g4175,
         g4176, g4177, g4178, g4179, g4180, g4181, g4191, g4192, g4193, g4194,
         g4195, g4196, g4197, g4198, g4199, g4200, g4201, g4202, g4203, g4204,
         g4205, g4206, g4207, g4208, g4209, g4210, g4211, g4212, g4213, g4214,
         g4215, g4216, g4887, g4888, g5101, g5105, g5658, g5659, g5816, g6253,
         g6254, g6255, g6256, g6257, g6258, g6259, g6260, g6261, g6262, g6263,
         g6264, g6265, g6266, g6267, g6268, g6269, g6270, g6271, g6272, g6273,
         g6274, g6275, g6276, g6277, g6278, g6279, g6280, g6281, g6282, g6283,
         g6284, g6285, g6842, g6920, g6926, g6932, g6942, g6949, g6955, g7744,
         g8061, g8062, g8271, g8313, g8316, g8318, g8323, g8328, g8331, g8335,
         g8340, g8347, g8349, g8352, g8561, g8562, g8563, g8564, g8565, g8566,
         g8976, g8977, g8978, g8979, g8980, g8981, g8982, g8983, g8984, g8985,
         g8986, g9451, g9961;
  wire   N599, g100, g101, g102, g103, g104, g1170, g1173, g1176, g1179, g1182,
         g1185, g1188, g1191, g1194, g1197, g1200, g1203, g18, g1960, g1961,
         g27, g28, g29, g30, g31, g41, g42, g43, g44, g45, g46, g47, g48, g82,
         g83, g84, g85, g86, g87, g872, g873, g88, g886, g889, g89, g892, g895,
         g898, g90, g901, g904, g907, g91, g910, g913, g916, g919, g92, g922,
         g925, g93, g94, g95, g96, g99, g1882, g312, g452, g11257, g123, g207,
         g713, g1558, g695, g461, g976, g709, g8432, g1092, g1574, g1864, g369,
         g1580, g39, g1424, g1672, g1077, g1231, g4, g774, g1304, g7290, g243,
         g1499, g1444, g757, g786, g1543, g315, g1534, g622, g1927, g1660,
         g278, g1436, g718, g8433, g554, g496, g11333, g981, g878, g590, g829,
         g1095, g704, g1265, g7302, g1786, g682, g8429, g1296, g7292, g587,
         g646, g327, g1389, g1371, g1956, g1955, g1675, g354, g639, g1684,
         g1791, g248, g1707, g351, g1604, g1098, g1896, g8282, g736, g8435,
         g1019, g1362, g745, g1419, g32, g876, g1086, g1486, g1730, g1504,
         g1470, g822, g583, g1678, g174, g1766, g1801, g186, g959, g1007,
         g1407, g1868, g758, g1718, g396, g11265, g1015, g38, g632, g1415,
         g1227, g1721, g16, g284, g426, g11256, g219, g806, g1428, g579, g1564,
         g225, g281, g1308, g611, g631, g1217, g1589, g1466, g1571, g1861,
         g1365, g1448, g1333, g153, g962, g766, g588, g486, g11331, g471,
         g1397, g580, g1950, g8288, g756, g755, g635, g549, g105, g1368, g1531,
         g1458, g572, g1011, g33, g1411, g1074, g444, g11259, g1474, g1080,
         g1713, g333, g269, g401, g11266, g1857, g9, g664, g965, g1400, g309,
         g814, g231, g557, g586, g869, g875, g1383, g158, g627, g1023, g259,
         g1361, g1206, g1327, g654, g293, g1346, g1633, g1508, g1240, g7297,
         g538, g11326, g416, g11269, g542, g11325, g1681, g374, g563, g1914,
         g8284, g530, g11328, g575, g1936, g1317, g1356, g357, g386, g11263,
         g1601, g166, g501, g11334, g262, g1840, g318, g794, g36, g302, g342,
         g1250, g7299, g1810, g1032, g1432, g1453, g363, g330, g35, g261, g516,
         g11337, g254, g778, g861, g1627, g1292, g7293, g290, g1850, g770,
         g1583, g466, g1561, g1546, g287, g560, g617, g17, g336, g456, g305,
         g345, g8, g1771, g865, g255, g1945, g1478, g1959, g1690, g1482, g296,
         g1663, g700, g8431, g360, g192, g1657, g722, g566, g1394, g1089,
         g1071, g986, g971, g143, g1814, g1212, g1918, g782, g1822, g237, g746,
         g1462, g178, g366, g837, g599, g1854, g944, g1941, g8287, g170, g1520,
         g686, g953, g1958, g40, g1733, g1270, g7303, g1796, g1324, g1540,
         g1377, g491, g11332, g1849, g213, g1781, g1900, g1245, g7298, g108,
         g630, g148, g833, g1923, g8285, g1314, g849, g1336, g272, g1806, g826,
         g1887, g8281, g37, g968, g1845, g1891, g1255, g7300, g257, g874, g591,
         g731, g636, g1218, g605, g182, g950, g857, g448, g11258, g1828, g1727,
         g1592, g1703, g1932, g8286, g1624, g1068, g578, g440, g11260, g476,
         g11338, g119, g668, g139, g34, g1848, g263, g818, g802, g275, g1524,
         g1577, g810, g391, g11264, g658, g1386, g253, g201, g1280, g7295,
         g1083, g650, g1636, g853, g421, g11270, g762, g956, g378, g589, g841,
         g1027, g1003, g1403, g1223, g406, g11267, g1811, g1654, g197, g1595,
         g1537, g727, g8434, g999, g798, g481, g11324, g754, g1330, g845, g790,
         g1490, g348, g868, g1260, g7301, g260, g131, g7, g258, g521, g11330,
         g1318, g1872, g677, g582, g1393, g1549, g947, g1834, g1598, g1321,
         g506, g11335, g546, g1909, g1552, g584, g1687, g1586, g324, g1341,
         g1710, g115, g135, g525, g11329, g581, g1607, g321, g1275, g11443,
         g1311, g1615, g382, g1374, g266, g1284, g7294, g1380, g673, g8428,
         g1853, g162, g411, g11268, g431, g11262, g1905, g8283, g1515, g1630,
         g991, g1300, g7291, g339, g256, g585, g1440, g1666, g1528, g1351,
         g127, g1618, g1235, g7296, g299, g435, g11261, g1555, g995, g1621,
         g643, g1494, g1567, g691, g8430, g534, g11327, g1776, g569, g1, g511,
         g11336, g1724, g12, g1878, g5529, g6551, g8054, g7709, g4940, g6481,
         g6215, g6529, g10707, g3435, g10408, g10336, g8940, g10855, g3399,
         g6907, g6155, g11647, g6910, g10417, g6828, g10800, g8019, g6821,
         g11478, g6516, g8244, g8631, g10793, g5910, g6824, g9931, g6759,
         g6502, g10797, g11625, g11372, g10771, g4114, g11293, g8173, g6533,
         g10405, g8245, g10767, g6000, g4903, g10720, g6934, g6123, g6838,
         g4905, g10798, g6830, g8944, g5543, g8921, g6096, g3431, g6733, g6823,
         g4890, g10863, g8039, g10664, g8923, g10712, g6755, g2791, g11514,
         g10411, g6902, g6015, g11340, g6542, g6507, g5556, g8505, g11641,
         g10765, g11305, g6126, g10414, g8060, g7191, g6469, g4893, g3418,
         g6901, g8043, g6929, g8049, g6786, g6234, g10864, g10862, g8051,
         g6541, g10773, g6523, g5404, g11393, g11561, g6908, g8768, g8885,
         g6333, g10515, g6045, g7590, g6468, g6672, g6840, g5914, g7705, g6038,
         g6471, g11303, g10663, g8920, g10788, g5396, g10583, g8045, g7843,
         g3425, g6537, g4902, g6080, g6059, g4089, g10866, g11603, g6332,
         g11488, g5918, g6894, g4076, g6534, g6928, g3414, g8055, g11291,
         g6833, g6918, g6915, g6911, g7441, g5996, g8047, g6832, g11481, g6478,
         g6897, g6042, g10402, g11609, g10859, g6054, g6508, g8050, g11376,
         g8559, g7032, g8767, g11483, g10776, g6513, g9272, g10898, g8052,
         g8766, g6205, g8820, g9124, g6839, g6522, g10936, g11320, g6841,
         g8769, g6224, g11349, g6470, g5755, g6515, g10791, g7632, g11485,
         g6331, g8053, g5763, g6480, g6795, g8938, g8775, g4891, g11290, g6501,
         g6334, g10719, g8765, g6916, g11308, g6820, g6922, g6747, g11391,
         g8649, g9555, g6071, g10858, g8926, g11602, g8041, g8922, g5536,
         g11605, g8048, g6528, g6524, g8046, g11482, g6923, g8937, g6538,
         g10339, g11306, g6895, g6163, g6179, g9721, g8776, g6827, g7244,
         g7586, g7930, g11300, g10718, g5445, g6088, g6679, g11636, g9266,
         g11608, g8059, g8771, g6035, g6198, g8973, g6834, g7134, g10795,
         g10770, g8773, g3462, g8939, g8772, g6093, g6500, g8777, g6244,
         g11640, g11487, g9110, g11380, g9269, g11314, g9150, g11298, g7202,
         g6819, g6243, g6514, g6983, g8040, g6900, g8042, g6546, g5770, g8889,
         g10711, g11312, g5287, g6479, g5849, g6656, g6906, g10717, g8770,
         g11610, g11604, g11486, g7581, g10799, g6439, g7133, g8044, g11607,
         g3506, g3407, g6193, g4904, g11292, g6822, g6912, g6898, g5421, g6924,
         g11310, g11294, g6026, g8024, g8945, g6525, g5083, g7541, g10860,
         g11579, g11639, g6826, g7626, g6829, g7660, g10722, g8887, g11484,
         g11286, g6002, g11606, g6757, g6216, g8941, g4892, g6930, g6049,
         g8943, g10861, g8779, g6180, g8774, g6099, g6831, g6068, g7137, g6545,
         g7257, g6909, g8384, g11392, g6506, g8883, g6728, g10724, n1005,
         n1007, n1008, n1010, n1012, n1013, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         g6955;
  assign g6280 = g100;
  assign g6281 = g101;
  assign g6282 = g102;
  assign g6283 = g103;
  assign g6284 = g104;
  assign g4205 = g1170;
  assign g4209 = g1173;
  assign g4210 = g1176;
  assign g4211 = g1179;
  assign g4212 = g1182;
  assign g4213 = g1185;
  assign g4214 = g1188;
  assign g4215 = g1191;
  assign g4216 = g1194;
  assign g4206 = g1197;
  assign g4207 = g1200;
  assign g4208 = g1203;
  assign g2355 = g18;
  assign g4888 = g1960;
  assign g4887 = g1961;
  assign g7744 = g27;
  assign g6285 = g28;
  assign g6253 = g29;
  assign g6254 = g30;
  assign g6255 = g31;
  assign g6256 = g41;
  assign g6257 = g42;
  assign g6258 = g43;
  assign g6259 = g44;
  assign g6260 = g45;
  assign g6261 = g46;
  assign g6262 = g47;
  assign g6263 = g48;
  assign g8335 = g82;
  assign g8328 = g82;
  assign g8349 = g82;
  assign g8352 = g82;
  assign g8313 = g82;
  assign g8318 = g82;
  assign g6264 = g82;
  assign g6265 = g83;
  assign g6266 = g84;
  assign g6267 = g85;
  assign g6268 = g86;
  assign g6269 = g87;
  assign g8061 = g872;
  assign g5101 = g872;
  assign g8062 = g873;
  assign g5105 = g873;
  assign g6270 = g88;
  assign g4191 = g886;
  assign g4192 = g889;
  assign g6271 = g89;
  assign g4193 = g892;
  assign g4194 = g895;
  assign g4195 = g898;
  assign g6272 = g90;
  assign g4197 = g901;
  assign g4198 = g904;
  assign g4199 = g907;
  assign g6273 = g91;
  assign g4200 = g910;
  assign g4201 = g913;
  assign g4202 = g916;
  assign g4203 = g919;
  assign g6274 = g92;
  assign g4204 = g922;
  assign g4196 = g925;
  assign g6275 = g93;
  assign g6276 = g94;
  assign g6277 = g95;
  assign g6278 = g96;
  assign g6279 = g99;
  assign g4177 = g774;
  assign g4180 = g786;
  assign g3007 = g878;
  assign g2602 = g587;
  assign g2609 = g583;
  assign g4173 = g758;
  assign g2605 = g579;
  assign g4175 = g766;
  assign g2603 = g588;
  assign g2606 = g580;
  assign g2612 = g586;
  assign g3069 = g1206;
  assign g5816 = g1810;
  assign g8271 = g1810;
  assign g4178 = g778;
  assign g4176 = g770;
  assign g2648 = g865;
  assign g4179 = g782;
  assign g2601 = g578;
  assign g4174 = g762;
  assign g2604 = g589;
  assign g4172 = g754;
  assign g4181 = g790;
  assign g2608 = g582;
  assign g2610 = g584;
  assign g2607 = g581;
  assign g2611 = g585;
  assign g8565 = g3435;
  assign g6949 = g3435;
  assign g10459 = g10408;
  assign g10377 = g10336;
  assign g8561 = g3399;
  assign g6920 = g3399;
  assign g10465 = g10417;
  assign g9961 = g9931;
  assign g9451 = g9931;
  assign g10457 = g10405;
  assign g8564 = g3431;
  assign g6942 = g3431;
  assign g10801 = g10712;
  assign g4171 = g2791;
  assign g10461 = g10411;
  assign g10463 = g10414;
  assign g5659 = g3418;
  assign g10628 = g10515;
  assign g11206 = g10583;
  assign g8563 = g3425;
  assign g6932 = g3425;
  assign g8562 = g3414;
  assign g6926 = g3414;
  assign g10455 = g10402;
  assign g10379 = g10339;
  assign g6842 = g5287;
  assign g5658 = g3407;
  assign g11489 = 1'b0;
  assign g8566 = g6955;
  assign g8981 = 1'b0;
  assign g8986 = 1'b0;
  assign g2986 = 1'b0;
  assign g8983 = 1'b0;
  assign g8979 = 1'b0;
  assign g8977 = 1'b0;
  assign g8985 = 1'b0;
  assign g8331 = 1'b1;
  assign g8347 = 1'b1;
  assign g8316 = 1'b1;
  assign g8340 = 1'b1;
  assign g8323 = 1'b1;
  assign g8984 = 1'b1;
  assign g8976 = 1'b1;
  assign g8982 = 1'b1;
  assign g8980 = 1'b1;
  assign g8978 = 1'b1;

  dff_533 DFF_1 ( .clk(CK), .q(g1882), .d(g8943) );
  dff_532 DFF_2 ( .clk(CK), .q(g312), .d(g255) );
  dff_531 DFF_3 ( .clk(CK), .q(g452), .d(g11257) );
  dff_530 DFF_4 ( .clk(CK), .q(g123), .d(g7032) );
  dff_529 DFF_5 ( .clk(CK), .q(g207), .d(g6830) );
  dff_528 DFF_6 ( .clk(CK), .q(g713), .d(g8920) );
  dff_524 DFF_10 ( .clk(CK), .q(g1558), .d(g6538) );
  dff_523 DFF_11 ( .clk(CK), .q(g695), .d(g8887) );
  dff_522 DFF_12 ( .clk(CK), .q(g461), .d(g11372) );
  dff_520 DFF_14 ( .clk(CK), .q(g976), .d(g11391) );
  dff_519 DFF_15 ( .clk(CK), .q(g709), .d(g8432) );
  dff_518 DFF_16 ( .clk(CK), .q(g1092), .d(g6088) );
  dff_517 DFF_17 ( .clk(CK), .q(g1574), .d(g6478) );
  dff_516 DFF_18 ( .clk(CK), .q(g1864), .d(g6795) );
  dff_515 DFF_19 ( .clk(CK), .q(g369), .d(g11320) );
  dff_514 DFF_20 ( .clk(CK), .q(g1580), .d(g6500) );
  dff_512 DFF_22 ( .clk(CK), .q(g39), .d_BAR(n1352) );
  dff_510 DFF_24 ( .clk(CK), .q(g1424), .d(g6216) );
  dff_508 DFF_26 ( .clk(CK), .q(g1672), .d(g10858) );
  dff_507 DFF_27 ( .clk(CK), .q(g1077), .d(g5914) );
  dff_506 DFF_28 ( .clk(CK), .q(g1231), .d(g7590) );
  dff_505 DFF_29 ( .clk(CK), .q(g4), .d(g6656) );
  dff_504 DFF_30 ( .clk(CK), .q(g774), .d(g6728) );
  dff_502 DFF_32 ( .clk(CK), .q(g1304), .d(g7290) );
  dff_501 DFF_33 ( .clk(CK), .q(g243), .d(g6841) );
  dff_500 DFF_34 ( .clk(CK), .q(g1499), .d(g8041) );
  dff_498 DFF_36 ( .clk(CK), .q(g1444), .d(g8766) );
  dff_497 DFF_37 ( .clk(CK), .q(g757), .d(g10788) );
  dff_496 DFF_38 ( .clk(CK), .q(g786), .d(g8019) );
  dff_495 DFF_39 ( .clk(CK), .q(g1543), .d(g6545) );
  dff_493 DFF_41 ( .clk(CK), .q(g315), .d(g256) );
  dff_492 DFF_42 ( .clk(CK), .q(g1534), .d(g6533) );
  dff_491 DFF_43 ( .clk(CK), .q(g622), .d(g8820) );
  dff_490 DFF_44 ( .clk(CK), .q(g1927), .d(g8941) );
  dff_489 DFF_45 ( .clk(CK), .q(g1660), .d(g10859) );
  dff_488 DFF_46 ( .clk(CK), .q(g278), .d(g6922) );
  dff_487 DFF_47 ( .clk(CK), .q(g1436), .d(g8772) );
  dff_486 DFF_48 ( .clk(CK), .q(g718), .d(g8433) );
  dff_484 DFF_50 ( .clk(CK), .q(g554), .d(g10793) );
  dff_483 DFF_51 ( .clk(CK), .q(g496), .d(g11333) );
  dff_482 DFF_52 ( .clk(CK), .q(g981), .d(g11392) );
  dff_481 DFF_53 ( .clk(CK), .q(g878), .d(g3506) );
  dff_480 DFF_54 ( .clk(CK), .q(g590), .d(g1713) );
  dff_479 DFF_55 ( .clk(CK), .q(g829), .d(g794) );
  dff_478 DFF_56 ( .clk(CK), .q(g1095), .d(g6093) );
  dff_477 DFF_57 ( .clk(CK), .q(g704), .d(g8889) );
  dff_476 DFF_58 ( .clk(CK), .q(g1265), .d(g7302) );
  dff_475 DFF_59 ( .clk(CK), .q(g1786), .d(g6525) );
  dff_474 DFF_60 ( .clk(CK), .q(g682), .d(g8429) );
  dff_473 DFF_61 ( .clk(CK), .q(g1296), .d(g7292) );
  dff_472 DFF_62 ( .clk(CK), .q(g587), .d(g104) );
  dff_470 DFF_64 ( .clk(CK), .q(g646), .d(g7134) );
  dff_469 DFF_65 ( .clk(CK), .q(g327), .d(g260) );
  dff_468 DFF_66 ( .clk(CK), .q(g1389), .d(g6333) );
  dff_467 DFF_67 ( .clk(CK), .q(g1371), .d(g6826) );
  dff_466 DFF_68 ( .clk(CK), .q(g1956), .d(g1955) );
  dff_465 DFF_69 ( .clk(CK), .q(g1675), .d(g10860) );
  dff_464 DFF_70 ( .clk(CK), .q(g354), .d(g11483) );
  dff_462 DFF_72 ( .clk(CK), .q(g639), .d(g7626) );
  dff_461 DFF_73 ( .clk(CK), .q(g1684), .d(g10866) );
  dff_459 DFF_75 ( .clk(CK), .q(g1791), .d(g6983) );
  dff_458 DFF_76 ( .clk(CK), .q(g248), .d(g6839) );
  dff_457 DFF_77 ( .clk(CK), .q(g1707), .d(g4076) );
  dff_455 DFF_79 ( .clk(CK), .q(g351), .d(g11482) );
  dff_454 DFF_80 ( .clk(CK), .q(g1957), .d(g1956) );
  dff_453 DFF_81 ( .clk(CK), .q(g1604), .d(g6507) );
  dff_452 DFF_82 ( .clk(CK), .q(g1098), .d(g6096) );
  dff_449 DFF_85 ( .clk(CK), .q(g1896), .d(g8282) );
  dff_448 DFF_86 ( .clk(CK), .q(g736), .d(g8435) );
  dff_447 DFF_87 ( .clk(CK), .q(g1019), .d(g6924) );
  dff_446 DFF_88 ( .clk(CK), .q(g1362), .d(g6819) );
  dff_445 DFF_89 ( .clk(CK), .q(g745), .d(g746) );
  dff_444 DFF_90 ( .clk(CK), .q(g1419), .d(g6244) );
  dff_442 DFF_92 ( .clk(CK), .q(g32), .d(g11286) );
  dff_441 DFF_93 ( .clk(CK), .d(g878), .q_BAR(g876) );
  dff_440 DFF_94 ( .clk(CK), .q(g1086), .d(g6071) );
  dff_439 DFF_95 ( .clk(CK), .q(g1486), .d(g8046) );
  dff_438 DFF_96 ( .clk(CK), .q(g1730), .d(g10707) );
  dff_437 DFF_97 ( .clk(CK), .q(g1504), .d(g6198) );
  dff_436 DFF_98 ( .clk(CK), .q(g1470), .d(g8051) );
  dff_435 DFF_99 ( .clk(CK), .q(g822), .d(g8024) );
  dff_434 DFF_100 ( .clk(CK), .q(g583), .d(g29) );
  dff_433 DFF_101 ( .clk(CK), .q(g1678), .d(g10862) );
  dff_432 DFF_102 ( .clk(CK), .q(g174), .d(g8050) );
  dff_431 DFF_103 ( .clk(CK), .q(g1766), .d(g7133) );
  dff_430 DFF_104 ( .clk(CK), .q(g1801), .d(g7930) );
  dff_429 DFF_105 ( .clk(CK), .q(g186), .d(g6832) );
  dff_428 DFF_106 ( .clk(CK), .q(g959), .d(g11308) );
  dff_426 DFF_108 ( .clk(CK), .q(g1007), .d(g6918) );
  dff_425 DFF_109 ( .clk(CK), .q(g1407), .d(g8769) );
  dff_423 DFF_111 ( .clk(CK), .q(g1868), .d(g6909) );
  dff_422 DFF_112 ( .clk(CK), .q(g758), .d(g4940) );
  dff_421 DFF_113 ( .clk(CK), .q(g1718), .d(g5404) );
  dff_420 DFF_114 ( .clk(CK), .q(g396), .d(g11265) );
  dff_419 DFF_115 ( .clk(CK), .q(g1015), .d(g6930) );
  dff_418 DFF_116 ( .clk(CK), .q(g38), .d(n2029) );
  dff_417 DFF_117 ( .clk(CK), .q(g632), .d(g4891) );
  dff_416 DFF_118 ( .clk(CK), .q(g1415), .d(g6224) );
  dff_415 DFF_119 ( .clk(CK), .q(g1227), .d(g7586) );
  dff_414 DFF_120 ( .clk(CK), .q(g1721), .d(g10770) );
  dff_412 DFF_122 ( .clk(CK), .q(g16), .d(n1007) );
  dff_411 DFF_123 ( .clk(CK), .q(g284), .d(g6934) );
  dff_410 DFF_124 ( .clk(CK), .q(g426), .d(g11256) );
  dff_409 DFF_125 ( .clk(CK), .q(g219), .d(g6824) );
  dff_407 DFF_127 ( .clk(CK), .q(g806), .d(g6126) );
  dff_406 DFF_128 ( .clk(CK), .q(g1428), .d(g8767) );
  dff_405 DFF_129 ( .clk(CK), .q(g579), .d(g102) );
  dff_404 DFF_130 ( .clk(CK), .q(g1564), .d(g6546) );
  dff_402 DFF_132 ( .clk(CK), .q(g225), .d(g6823) );
  dff_401 DFF_133 ( .clk(CK), .q(g281), .d(g6928) );
  dff_400 DFF_134 ( .clk(CK), .q(g1308), .d(g11602) );
  dff_399 DFF_135 ( .clk(CK), .q(g611), .d(g9721) );
  dff_398 DFF_136 ( .clk(CK), .q(g631), .d(g4890) );
  dff_397 DFF_137 ( .clk(CK), .q(g1217), .d(n1010) );
  dff_396 DFF_138 ( .clk(CK), .q(g1589), .d(g6524) );
  dff_395 DFF_139 ( .clk(CK), .q(g1466), .d(g8045) );
  dff_394 DFF_140 ( .clk(CK), .q(g1571), .d(g6469) );
  dff_393 DFF_141 ( .clk(CK), .q(g1861), .d(g6471) );
  dff_392 DFF_142 ( .clk(CK), .q(g1365), .d(g6821) );
  dff_391 DFF_143 ( .clk(CK), .q(g1448), .d(g11514) );
  dff_388 DFF_146 ( .clk(CK), .q(g1333), .d(g11610) );
  dff_387 DFF_147 ( .clk(CK), .q(g153), .d(g7843) );
  dff_386 DFF_148 ( .clk(CK), .q(g962), .d(g11310) );
  dff_385 DFF_149 ( .clk(CK), .q(g766), .d(g5536) );
  dff_384 DFF_150 ( .clk(CK), .q(g588), .d(g28) );
  dff_383 DFF_151 ( .clk(CK), .q(g486), .d(g11331) );
  dff_382 DFF_152 ( .clk(CK), .q(g471), .d(g11380) );
  dff_381 DFF_153 ( .clk(CK), .q(g1397), .d(g6838) );
  dff_380 DFF_154 ( .clk(CK), .q(g580), .d(g103) );
  dff_379 DFF_155 ( .clk(CK), .q(g1950), .d(g8288) );
  dff_378 DFF_156 ( .clk(CK), .q(g756), .d(g755) );
  dff_377 DFF_157 ( .clk(CK), .q(g635), .d(g4892) );
  dff_375 DFF_159 ( .clk(CK), .q(g549), .d(g10855) );
  dff_373 DFF_161 ( .clk(CK), .q(g105), .d(g10898) );
  dff_371 DFF_163 ( .clk(CK), .q(g1368), .d(g6822) );
  dff_370 DFF_164 ( .clk(CK), .q(g1531), .d(g6528) );
  dff_369 DFF_165 ( .clk(CK), .q(g1458), .d(g6180) );
  dff_368 DFF_166 ( .clk(CK), .q(g572), .d(g10718) );
  dff_367 DFF_167 ( .clk(CK), .q(g1011), .d(g6912) );
  dff_366 DFF_168 ( .clk(CK), .q(g33), .d(g10719) );
  dff_365 DFF_169 ( .clk(CK), .q(g1411), .d(g6234) );
  dff_364 DFF_170 ( .clk(CK), .q(g1074), .d(g6099) );
  dff_363 DFF_171 ( .clk(CK), .q(g444), .d(g11259) );
  dff_362 DFF_172 ( .clk(CK), .q(g1474), .d(g8039) );
  dff_361 DFF_173 ( .clk(CK), .q(g1080), .d(g6059) );
  dff_360 DFF_174 ( .clk(CK), .q(g1713), .d(g5396) );
  dff_359 DFF_175 ( .clk(CK), .q(g333), .d(g262) );
  dff_358 DFF_176 ( .clk(CK), .q(g269), .d(g6906) );
  dff_357 DFF_177 ( .clk(CK), .q(g401), .d(g11266) );
  dff_356 DFF_178 ( .clk(CK), .q(g1857), .d(g11294) );
  dff_355 DFF_179 ( .clk(CK), .q(g9), .d(g5421) );
  dff_354 DFF_180 ( .clk(CK), .q(g664), .d(g8649) );
  dff_353 DFF_181 ( .clk(CK), .q(g965), .d(g11312) );
  dff_352 DFF_182 ( .clk(CK), .q(g1400), .d(g6840) );
  dff_351 DFF_183 ( .clk(CK), .q(g309), .d(g254) );
  dff_350 DFF_184 ( .clk(CK), .q(g814), .d(g7202) );
  dff_349 DFF_185 ( .clk(CK), .q(g231), .d(g6834) );
  dff_348 DFF_186 ( .clk(CK), .q(g557), .d(g10795) );
  dff_347 DFF_187 ( .clk(CK), .q(g586), .d(g103) );
  dff_346 DFF_188 ( .clk(CK), .q(g869), .d(g875) );
  dff_345 DFF_189 ( .clk(CK), .q(g1383), .d(g6831) );
  dff_344 DFF_190 ( .clk(CK), .q(g158), .d(g8060) );
  dff_343 DFF_191 ( .clk(CK), .q(g627), .d(g4893) );
  dff_342 DFF_192 ( .clk(CK), .q(g1023), .d(g7244) );
  dff_341 DFF_193 ( .clk(CK), .q(g259), .d(g6026) );
  dff_340 DFF_194 ( .clk(CK), .d(g1206), .q_BAR(g1361) );
  dff_339 DFF_195 ( .clk(CK), .q(g1327), .d(g11608) );
  dff_338 DFF_196 ( .clk(CK), .q(g654), .d(g7660) );
  dff_337 DFF_197 ( .clk(CK), .q(g293), .d(g6911) );
  dff_336 DFF_198 ( .clk(CK), .q(g1346), .d(g11640) );
  dff_335 DFF_199 ( .clk(CK), .q(g1633), .d(g8777) );
  dff_333 DFF_201 ( .clk(CK), .q(g1508), .d(g6215) );
  dff_332 DFF_202 ( .clk(CK), .q(g1240), .d(g7297) );
  dff_331 DFF_203 ( .clk(CK), .q(g538), .d(g11326) );
  dff_330 DFF_204 ( .clk(CK), .q(g416), .d(g11269) );
  dff_329 DFF_205 ( .clk(CK), .q(g542), .d(g11325) );
  dff_328 DFF_206 ( .clk(CK), .q(g1681), .d(g10864) );
  dff_327 DFF_207 ( .clk(CK), .q(g374), .d(g11290) );
  dff_326 DFF_208 ( .clk(CK), .q(g563), .d(g10798) );
  dff_325 DFF_209 ( .clk(CK), .q(g1914), .d(g8284) );
  dff_324 DFF_210 ( .clk(CK), .q(g530), .d(g11328) );
  dff_323 DFF_211 ( .clk(CK), .q(g575), .d(g10800) );
  dff_322 DFF_212 ( .clk(CK), .q(g1936), .d(g8944) );
  dff_319 DFF_215 ( .clk(CK), .d(g1356), .q_BAR(g1317) );
  dff_318 DFF_216 ( .clk(CK), .q(g357), .d(g11484) );
  dff_317 DFF_217 ( .clk(CK), .q(g386), .d(g11263) );
  dff_316 DFF_218 ( .clk(CK), .q(g1601), .d(g6501) );
  dff_314 DFF_220 ( .clk(CK), .q(g166), .d(g6757) );
  dff_313 DFF_221 ( .clk(CK), .q(g501), .d(g11334) );
  dff_312 DFF_222 ( .clk(CK), .q(g262), .d(g6042) );
  dff_311 DFF_223 ( .clk(CK), .q(g1840), .d(g8384) );
  dff_309 DFF_225 ( .clk(CK), .q(g318), .d(g257) );
  dff_308 DFF_226 ( .clk(CK), .q(g1356), .d(g5763) );
  dff_307 DFF_227 ( .clk(CK), .q(g794), .d(g5849) );
  dff_306 DFF_228 ( .clk(CK), .q(g36), .d_BAR(n1341) );
  dff_305 DFF_229 ( .clk(CK), .q(g302), .d(g6929) );
  dff_304 DFF_230 ( .clk(CK), .q(g342), .d(g11488) );
  dff_303 DFF_231 ( .clk(CK), .q(g1250), .d(g7299) );
  dff_301 DFF_233 ( .clk(CK), .d(g1958), .q_BAR(g1810) );
  dff_300 DFF_234 ( .clk(CK), .q(g1032), .d(g7257) );
  dff_299 DFF_235 ( .clk(CK), .q(g1432), .d(g8775) );
  dff_297 DFF_237 ( .clk(CK), .q(g1453), .d(g5770) );
  dff_296 DFF_238 ( .clk(CK), .q(g363), .d(g11486) );
  dff_295 DFF_239 ( .clk(CK), .q(g330), .d(g261) );
  dff_292 DFF_242 ( .clk(CK), .q(g35), .d(n1354) );
  dff_290 DFF_244 ( .clk(CK), .q(g261), .d(g6038) );
  dff_289 DFF_245 ( .clk(CK), .q(g516), .d(g11337) );
  dff_288 DFF_246 ( .clk(CK), .q(g254), .d(g6045) );
  dff_287 DFF_247 ( .clk(CK), .q(g778), .d(g7191) );
  dff_286 DFF_248 ( .clk(CK), .q(g861), .d(g826) );
  dff_285 DFF_249 ( .clk(CK), .d(g8774), .q_BAR(g1627) );
  dff_284 DFF_250 ( .clk(CK), .q(g1292), .d(g7293) );
  dff_283 DFF_251 ( .clk(CK), .q(g290), .d(g6907) );
  dff_282 DFF_252 ( .clk(CK), .q(g1850), .d(g4903) );
  dff_281 DFF_253 ( .clk(CK), .q(g770), .d(g6123) );
  dff_280 DFF_254 ( .clk(CK), .q(g1583), .d(g6506) );
  dff_279 DFF_255 ( .clk(CK), .q(g466), .d(g11376) );
  dff_278 DFF_256 ( .clk(CK), .q(g1561), .d(g6542) );
  dff_276 DFF_258 ( .clk(CK), .q(g1546), .d(g6551) );
  dff_275 DFF_259 ( .clk(CK), .q(g287), .d(g6901) );
  dff_274 DFF_260 ( .clk(CK), .q(g560), .d(g10797) );
  dff_273 DFF_261 ( .clk(CK), .q(g617), .d(g8505) );
  dff_272 DFF_262 ( .clk(CK), .q(g17), .d(n1005) );
  dff_271 DFF_263 ( .clk(CK), .q(g336), .d(g11647) );
  dff_270 DFF_264 ( .clk(CK), .q(g456), .d(g11340) );
  dff_269 DFF_265 ( .clk(CK), .d(g253), .q_BAR(g305) );
  dff_268 DFF_266 ( .clk(CK), .q(g345), .d(g11625) );
  dff_267 DFF_267 ( .clk(CK), .q(g8), .d(g636) );
  dff_266 DFF_268 ( .clk(CK), .q(g1771), .d(g6502) );
  dff_265 DFF_269 ( .clk(CK), .q(g865), .d(N599) );
  dff_264 DFF_270 ( .clk(CK), .q(g255), .d(g6049) );
  dff_263 DFF_271 ( .clk(CK), .q(g1945), .d(g8945) );
  dff_261 DFF_273 ( .clk(CK), .q(g1478), .d(g8040) );
  dff_259 DFF_275 ( .clk(CK), .q(g1959), .d(n1008) );
  dff_258 DFF_276 ( .clk(CK), .q(g1690), .d(g6155) );
  dff_257 DFF_277 ( .clk(CK), .q(g1482), .d(g8043) );
  dff_255 DFF_279 ( .clk(CK), .q(g296), .d(g6916) );
  dff_254 DFF_280 ( .clk(CK), .q(g1663), .d(g10861) );
  dff_253 DFF_281 ( .clk(CK), .q(g700), .d(g8431) );
  dff_251 DFF_283 ( .clk(CK), .q(g360), .d(g11485) );
  dff_250 DFF_284 ( .clk(CK), .q(g192), .d(g6334) );
  dff_249 DFF_285 ( .clk(CK), .q(g1657), .d(g10767) );
  dff_248 DFF_286 ( .clk(CK), .q(g722), .d(g8923) );
  dff_246 DFF_288 ( .clk(CK), .q(g566), .d(g10799) );
  dff_245 DFF_289 ( .clk(CK), .q(g1394), .d(g6747) );
  dff_244 DFF_290 ( .clk(CK), .q(g1089), .d(g6080) );
  dff_242 DFF_292 ( .clk(CK), .q(g1071), .d(g5910) );
  dff_241 DFF_293 ( .clk(CK), .q(g986), .d(g11393) );
  dff_240 DFF_294 ( .clk(CK), .q(g971), .d(g11349) );
  dff_239 DFF_295 ( .clk(CK), .q(g1955), .d(g83) );
  dff_238 DFF_296 ( .clk(CK), .q(g143), .d(g6439) );
  dff_237 DFF_297 ( .clk(CK), .q(g1814), .d(g9266) );
  dff_235 DFF_299 ( .clk(CK), .q(g1212), .d(g1217) );
  dff_234 DFF_300 ( .clk(CK), .q(g1918), .d(g8940) );
  dff_233 DFF_301 ( .clk(CK), .q(g782), .d(g7705) );
  dff_232 DFF_302 ( .clk(CK), .q(g1822), .d(g9269) );
  dff_231 DFF_303 ( .clk(CK), .q(g237), .d(g6820) );
  dff_230 DFF_304 ( .clk(CK), .q(g746), .d(g756) );
  dff_228 DFF_306 ( .clk(CK), .q(g1462), .d(g8042) );
  dff_227 DFF_307 ( .clk(CK), .q(g178), .d(g6759) );
  dff_226 DFF_308 ( .clk(CK), .q(g366), .d(g11487) );
  dff_225 DFF_309 ( .clk(CK), .q(g837), .d(g802) );
  dff_224 DFF_310 ( .clk(CK), .q(g599), .d(g9124) );
  dff_223 DFF_311 ( .clk(CK), .q(g1854), .d(g11293) );
  dff_222 DFF_312 ( .clk(CK), .q(g944), .d(g11298) );
  dff_221 DFF_313 ( .clk(CK), .q(g1941), .d(g8287) );
  dff_220 DFF_314 ( .clk(CK), .q(g170), .d(g8047) );
  dff_219 DFF_315 ( .clk(CK), .q(g1520), .d(g6205) );
  dff_218 DFF_316 ( .clk(CK), .q(g686), .d(g8885) );
  dff_217 DFF_317 ( .clk(CK), .q(g953), .d(g11305) );
  dff_216 DFF_318 ( .clk(CK), .q(g1958), .d(g5556) );
  dff_215 DFF_319 ( .clk(CK), .q(g40), .d(g10664) );
  dff_213 DFF_321 ( .clk(CK), .q(g1733), .d(g10711) );
  dff_212 DFF_322 ( .clk(CK), .q(g1270), .d(g7303) );
  dff_210 DFF_324 ( .clk(CK), .q(g1796), .d(g7541) );
  dff_209 DFF_325 ( .clk(CK), .q(g1324), .d(g11607) );
  dff_208 DFF_326 ( .clk(CK), .q(g1540), .d(g6541) );
  dff_207 DFF_327 ( .clk(CK), .q(g1377), .d(g6827) );
  dff_206 DFF_328 ( .clk(CK), .q(g1206), .d(g4114) );
  dff_205 DFF_329 ( .clk(CK), .q(g491), .d(g11332) );
  dff_204 DFF_330 ( .clk(CK), .q(g1849), .d(g4902) );
  dff_203 DFF_331 ( .clk(CK), .q(g213), .d(g6828) );
  dff_202 DFF_332 ( .clk(CK), .q(g1781), .d(g6516) );
  dff_201 DFF_333 ( .clk(CK), .q(g1900), .d(g8938) );
  dff_200 DFF_334 ( .clk(CK), .q(g1245), .d(g7298) );
  dff_199 DFF_335 ( .clk(CK), .q(g108), .d(g11561) );
  dff_198 DFF_336 ( .clk(CK), .q(g630), .d(g6672) );
  dff_197 DFF_337 ( .clk(CK), .q(g148), .d(g8048) );
  dff_196 DFF_338 ( .clk(CK), .q(g833), .d(g798) );
  dff_195 DFF_339 ( .clk(CK), .q(g1923), .d(g8285) );
  dff_192 DFF_342 ( .clk(CK), .q(g1314), .d(g11604) );
  dff_191 DFF_343 ( .clk(CK), .q(g849), .d(g814) );
  dff_190 DFF_344 ( .clk(CK), .q(g1336), .d(g11636) );
  dff_189 DFF_345 ( .clk(CK), .q(g272), .d(g6910) );
  dff_188 DFF_346 ( .clk(CK), .q(g1806), .d(g8173) );
  dff_187 DFF_347 ( .clk(CK), .q(g826), .d(g8245) );
  dff_185 DFF_349 ( .clk(CK), .q(g1887), .d(g8281) );
  dff_184 DFF_350 ( .clk(CK), .q(g37), .d_BAR(n1342) );
  dff_183 DFF_351 ( .clk(CK), .q(g968), .d(g11314) );
  dff_182 DFF_352 ( .clk(CK), .q(g1845), .d(g4905) );
  dff_180 DFF_354 ( .clk(CK), .q(g1891), .d(g8937) );
  dff_179 DFF_355 ( .clk(CK), .q(g1255), .d(g7300) );
  dff_178 DFF_356 ( .clk(CK), .q(g257), .d(g6002) );
  dff_177 DFF_357 ( .clk(CK), .q(g874), .d(n1012) );
  dff_176 DFF_358 ( .clk(CK), .q(g591), .d(g9110) );
  dff_175 DFF_359 ( .clk(CK), .q(g731), .d(g8926) );
  dff_174 DFF_360 ( .clk(CK), .q(g636), .d(g8631) );
  dff_173 DFF_361 ( .clk(CK), .q(g1218), .d(g7632) );
  dff_172 DFF_362 ( .clk(CK), .q(g605), .d(g9150) );
  dff_170 DFF_364 ( .clk(CK), .q(g182), .d(g6786) );
  dff_169 DFF_365 ( .clk(CK), .q(g950), .d(g11303) );
  dff_167 DFF_367 ( .clk(CK), .q(g857), .d(g822) );
  dff_166 DFF_368 ( .clk(CK), .q(g448), .d(g11258) );
  dff_165 DFF_369 ( .clk(CK), .q(g1828), .d(g9272) );
  dff_164 DFF_370 ( .clk(CK), .q(g1727), .d(g10773) );
  dff_163 DFF_371 ( .clk(CK), .q(g1592), .d(g6470) );
  dff_162 DFF_372 ( .clk(CK), .q(g1703), .d(g5083) );
  dff_161 DFF_373 ( .clk(CK), .q(g1932), .d(g8286) );
  dff_160 DFF_374 ( .clk(CK), .d(g8773), .q_BAR(g1624) );
  dff_158 DFF_376 ( .clk(CK), .q(g1068), .d(g6054) );
  dff_157 DFF_377 ( .clk(CK), .q(g578), .d(g101) );
  dff_156 DFF_378 ( .clk(CK), .q(g440), .d(g11260) );
  dff_155 DFF_379 ( .clk(CK), .q(g476), .d(g11338) );
  dff_154 DFF_380 ( .clk(CK), .q(g119), .d(g5918) );
  dff_153 DFF_381 ( .clk(CK), .q(g668), .d(g8922) );
  dff_152 DFF_382 ( .clk(CK), .q(g139), .d(g8049) );
  dff_150 DFF_384 ( .clk(CK), .q(g34), .d(g10720) );
  dff_149 DFF_385 ( .clk(CK), .q(g1848), .d(g6755) );
  dff_148 DFF_386 ( .clk(CK), .q(g263), .d(g6897) );
  dff_147 DFF_387 ( .clk(CK), .q(g818), .d(g7709) );
  dff_145 DFF_389 ( .clk(CK), .q(g802), .d(g5543) );
  dff_144 DFF_390 ( .clk(CK), .q(g275), .d(g6915) );
  dff_143 DFF_391 ( .clk(CK), .q(g1524), .d(g6513) );
  dff_142 DFF_392 ( .clk(CK), .q(g1577), .d(g6480) );
  dff_141 DFF_393 ( .clk(CK), .q(g810), .d(g6733) );
  dff_140 DFF_394 ( .clk(CK), .q(g391), .d(g11264) );
  dff_139 DFF_395 ( .clk(CK), .q(g658), .d(g8973) );
  dff_138 DFF_396 ( .clk(CK), .q(g1386), .d(g6833) );
  dff_137 DFF_397 ( .clk(CK), .q(g253), .d(g5996) );
  dff_136 DFF_398 ( .clk(CK), .q(g875), .d(n1013) );
  dff_134 DFF_400 ( .clk(CK), .d(g5755), .q_BAR(g201) );
  dff_133 DFF_401 ( .clk(CK), .q(g1280), .d(g7295) );
  dff_132 DFF_402 ( .clk(CK), .q(g1083), .d(g6068) );
  dff_131 DFF_403 ( .clk(CK), .q(g650), .d(g7137) );
  dff_130 DFF_404 ( .clk(CK), .q(g1636), .d(g8779) );
  dff_129 DFF_405 ( .clk(CK), .q(g853), .d(g818) );
  dff_128 DFF_406 ( .clk(CK), .q(g421), .d(g11270) );
  dff_127 DFF_407 ( .clk(CK), .q(g762), .d(g5529) );
  dff_126 DFF_408 ( .clk(CK), .q(g956), .d(g11306) );
  dff_125 DFF_409 ( .clk(CK), .q(g378), .d(g11291) );
  dff_123 DFF_411 ( .clk(CK), .q(g589), .d(g29) );
  dff_122 DFF_412 ( .clk(CK), .q(g841), .d(g806) );
  dff_121 DFF_413 ( .clk(CK), .q(g1027), .d(g6894) );
  dff_120 DFF_414 ( .clk(CK), .q(g1003), .d(g6902) );
  dff_119 DFF_415 ( .clk(CK), .q(g1403), .d(g8765) );
  dff_116 DFF_418 ( .clk(CK), .q(g1223), .d(g7581) );
  dff_115 DFF_419 ( .clk(CK), .q(g406), .d(g11267) );
  dff_114 DFF_420 ( .clk(CK), .q(g1811), .d(g10936) );
  dff_111 DFF_423 ( .clk(CK), .q(g1654), .d(g10765) );
  dff_110 DFF_424 ( .clk(CK), .q(g197), .d(g6332) );
  dff_109 DFF_425 ( .clk(CK), .q(g1595), .d(g6479) );
  dff_108 DFF_426 ( .clk(CK), .q(g1537), .d(g6537) );
  dff_107 DFF_427 ( .clk(CK), .q(g727), .d(g8434) );
  dff_106 DFF_428 ( .clk(CK), .q(g999), .d(g6908) );
  dff_105 DFF_429 ( .clk(CK), .q(g798), .d(g6243) );
  dff_104 DFF_430 ( .clk(CK), .q(g481), .d(g11324) );
  dff_103 DFF_431 ( .clk(CK), .q(g754), .d(g3462) );
  dff_102 DFF_432 ( .clk(CK), .q(g1330), .d(g11609) );
  dff_101 DFF_433 ( .clk(CK), .q(g845), .d(g810) );
  dff_100 DFF_434 ( .clk(CK), .q(g790), .d(g8244) );
  dff_97 DFF_437 ( .clk(CK), .q(g1490), .d(g8052) );
  dff_94 DFF_440 ( .clk(CK), .q(g348), .d(g11481) );
  dff_93 DFF_441 ( .clk(CK), .q(g868), .d(g874) );
  dff_92 DFF_442 ( .clk(CK), .q(g1260), .d(g7301) );
  dff_91 DFF_443 ( .clk(CK), .q(g260), .d(g6035) );
  dff_90 DFF_444 ( .clk(CK), .q(g131), .d(g8059) );
  dff_89 DFF_445 ( .clk(CK), .q(g7), .d(g1854) );
  dff_88 DFF_446 ( .clk(CK), .q(g258), .d(g6015) );
  dff_87 DFF_447 ( .clk(CK), .q(g521), .d(g11330) );
  dff_86 DFF_448 ( .clk(CK), .q(g1318), .d(g11605) );
  dff_85 DFF_449 ( .clk(CK), .q(g1872), .d(g8921) );
  dff_84 DFF_450 ( .clk(CK), .q(g677), .d(g8883) );
  dff_83 DFF_451 ( .clk(CK), .q(g582), .d(g28) );
  dff_82 DFF_452 ( .clk(CK), .q(g1393), .d(g6163) );
  dff_81 DFF_453 ( .clk(CK), .q(g1549), .d(g6523) );
  dff_80 DFF_454 ( .clk(CK), .q(g947), .d(g11300) );
  dff_79 DFF_455 ( .clk(CK), .q(g1834), .d(g9555) );
  dff_78 DFF_456 ( .clk(CK), .q(g1598), .d(g6481) );
  dff_76 DFF_458 ( .clk(CK), .q(g1321), .d(g11606) );
  dff_75 DFF_459 ( .clk(CK), .q(g506), .d(g11335) );
  dff_74 DFF_460 ( .clk(CK), .q(g546), .d(g10791) );
  dff_73 DFF_461 ( .clk(CK), .q(g1909), .d(g8939) );
  dff_72 DFF_462 ( .clk(CK), .q(g755), .d(g83) );
  dff_71 DFF_463 ( .clk(CK), .q(g1552), .d(g6529) );
  dff_70 DFF_464 ( .clk(CK), .q(g584), .d(g101) );
  dff_69 DFF_465 ( .clk(CK), .q(g1687), .d(g10776) );
  dff_68 DFF_466 ( .clk(CK), .q(g1586), .d(g6514) );
  dff_67 DFF_467 ( .clk(CK), .q(g324), .d(g259) );
  dff_64 DFF_470 ( .clk(CK), .q(g1341), .d(g11639) );
  dff_63 DFF_471 ( .clk(CK), .q(g1710), .d(g4089) );
  dff_61 DFF_473 ( .clk(CK), .q(g115), .d(g6179) );
  dff_60 DFF_474 ( .clk(CK), .q(g135), .d(g8053) );
  dff_59 DFF_475 ( .clk(CK), .q(g525), .d(g11329) );
  dff_58 DFF_476 ( .clk(CK), .q(g581), .d(g104) );
  dff_57 DFF_477 ( .clk(CK), .q(g1607), .d(g6515) );
  dff_56 DFF_478 ( .clk(CK), .q(g321), .d(g258) );
  dff_54 DFF_480 ( .clk(CK), .q(g1275), .d(g11443) );
  dff_53 DFF_481 ( .clk(CK), .q(g1311), .d(g11603) );
  dff_52 DFF_482 ( .clk(CK), .d(g8770), .q_BAR(g1615) );
  dff_51 DFF_483 ( .clk(CK), .q(g382), .d(g11292) );
  dff_50 DFF_484 ( .clk(CK), .q(g1374), .d(g6331) );
  dff_49 DFF_485 ( .clk(CK), .q(g266), .d(g6900) );
  dff_48 DFF_486 ( .clk(CK), .q(g1284), .d(g7294) );
  dff_47 DFF_487 ( .clk(CK), .q(g1380), .d(g6829) );
  dff_46 DFF_488 ( .clk(CK), .q(g673), .d(g8428) );
  dff_45 DFF_489 ( .clk(CK), .q(g1853), .d(g4904) );
  dff_44 DFF_490 ( .clk(CK), .q(g162), .d(g8054) );
  dff_43 DFF_491 ( .clk(CK), .q(g411), .d(g11268) );
  dff_42 DFF_492 ( .clk(CK), .q(g431), .d(g11262) );
  dff_41 DFF_493 ( .clk(CK), .q(g1905), .d(g8283) );
  dff_40 DFF_494 ( .clk(CK), .q(g1515), .d(g6193) );
  dff_39 DFF_495 ( .clk(CK), .q(g1630), .d(g8776) );
  dff_37 DFF_497 ( .clk(CK), .q(g991), .d(g6898) );
  dff_36 DFF_498 ( .clk(CK), .q(g1300), .d(g7291) );
  dff_35 DFF_499 ( .clk(CK), .q(g339), .d(g11478) );
  dff_34 DFF_500 ( .clk(CK), .q(g256), .d(g6000) );
  dff_32 DFF_502 ( .clk(CK), .q(g585), .d(g102) );
  dff_31 DFF_503 ( .clk(CK), .q(g1440), .d(g8768) );
  dff_30 DFF_504 ( .clk(CK), .q(g1666), .d(g10863) );
  dff_29 DFF_505 ( .clk(CK), .q(g1528), .d(g6522) );
  dff_28 DFF_506 ( .clk(CK), .q(g1351), .d(g11641) );
  dff_26 DFF_508 ( .clk(CK), .q(g127), .d(g8044) );
  dff_25 DFF_509 ( .clk(CK), .q(g1618), .d(g11579) );
  dff_24 DFF_510 ( .clk(CK), .q(g1235), .d(g7296) );
  dff_23 DFF_511 ( .clk(CK), .q(g299), .d(g6923) );
  dff_22 DFF_512 ( .clk(CK), .q(g435), .d(g11261) );
  dff_20 DFF_514 ( .clk(CK), .q(g1555), .d(g6534) );
  dff_19 DFF_515 ( .clk(CK), .q(g995), .d(g6895) );
  dff_18 DFF_516 ( .clk(CK), .q(g1621), .d(g8771) );
  dff_16 DFF_518 ( .clk(CK), .d(g7441), .q_BAR(g643) );
  dff_15 DFF_519 ( .clk(CK), .q(g1494), .d(g8055) );
  dff_14 DFF_520 ( .clk(CK), .q(g1567), .d(g6468) );
  dff_13 DFF_521 ( .clk(CK), .q(g691), .d(g8430) );
  dff_12 DFF_522 ( .clk(CK), .q(g534), .d(g11327) );
  dff_11 DFF_523 ( .clk(CK), .q(g1776), .d(g6508) );
  dff_10 DFF_524 ( .clk(CK), .q(g569), .d(g10717) );
  dff_6 DFF_528 ( .clk(CK), .q(g1), .d(g6679) );
  dff_5 DFF_529 ( .clk(CK), .q(g511), .d(g11336) );
  dff_4 DFF_530 ( .clk(CK), .q(g1724), .d(g10771) );
  dff_3 DFF_531 ( .clk(CK), .q(g12), .d(g5445) );
  dff_2 DFF_532 ( .clk(CK), .q(g1878), .d(g8559) );
  INVX0 U1518 ( .INP(n1467), .ZN(n1470) );
  NAND3X0 U1519 ( .IN1(g369), .IN2(n1250), .IN3(n1459), .QN(n1483) );
  AND2X1 U1520 ( .IN1(n1257), .IN2(n1256), .Q(n1026) );
  NAND2X1 U1521 ( .IN1(g10722), .IN2(g109), .QN(n1876) );
  INVX2 U1522 ( .INP(n1071), .ZN(n1207) );
  NAND3X0 U1523 ( .IN1(g971), .IN2(n1609), .IN3(g10788), .QN(n1586) );
  MUX21X1 U1524 ( .IN1(n1239), .IN2(g312), .S(n1245), .Q(n1769) );
  AND2X1 U1525 ( .IN1(g1546), .IN2(n1206), .Q(n1015) );
  XOR2X2 U1526 ( .IN1(n1264), .IN2(n1016), .Q(n1266) );
  MUX21X1 U1527 ( .IN1(g401), .IN2(g406), .S(n1968), .Q(g11267) );
  MUX21X1 U1528 ( .IN1(g396), .IN2(g401), .S(n1470), .Q(g11266) );
  NOR2X0 U1529 ( .IN1(g1703), .IN2(g1696), .QN(n2007) );
  MUX21X1 U1530 ( .IN1(n1981), .IN2(n1980), .S(n1470), .Q(n1982) );
  MUX21X1 U1531 ( .IN1(g448), .IN2(g444), .S(n1470), .Q(g11259) );
  MUX21X1 U1532 ( .IN1(g481), .IN2(g486), .S(n1470), .Q(g11331) );
  MUX21X1 U1533 ( .IN1(g444), .IN2(g440), .S(n1470), .Q(g11260) );
  OR3X1 U1534 ( .IN1(n1471), .IN2(n1470), .IN3(n1469), .Q(n1511) );
  MUX21X1 U1535 ( .IN1(g486), .IN2(g491), .S(n1470), .Q(g11332) );
  MUX21X1 U1536 ( .IN1(g435), .IN2(g431), .S(n1470), .Q(g11262) );
  MUX21X1 U1537 ( .IN1(g440), .IN2(g435), .S(n1470), .Q(g11261) );
  NAND2X0 U1538 ( .IN1(n1115), .IN2(n1129), .QN(g10719) );
  OAI22X1 U1539 ( .IN1(n1876), .IN2(n1744), .IN3(n1021), .IN4(n1743), .QN(
        n1424) );
  AND2X1 U1540 ( .IN1(n1354), .IN2(g10722), .Q(n1897) );
  AND3X1 U1541 ( .IN1(n1114), .IN2(n1113), .IN3(n1112), .Q(n1115) );
  AND4X1 U1542 ( .IN1(n1178), .IN2(n1177), .IN3(n1176), .IN4(n1193), .Q(n1179)
         );
  NAND3X0 U1543 ( .IN1(n1349), .IN2(n1348), .IN3(n1347), .QN(n1350) );
  NAND4X0 U1544 ( .IN1(n1346), .IN2(n1345), .IN3(n1344), .IN4(n1343), .QN(
        n1351) );
  AND2X1 U1545 ( .IN1(n1304), .IN2(g1327), .Q(n1305) );
  AND2X1 U1546 ( .IN1(n1832), .IN2(n1273), .Q(n1274) );
  NAND3X0 U1547 ( .IN1(n1739), .IN2(g1828), .IN3(n1798), .QN(n1740) );
  AND2X1 U1548 ( .IN1(n2008), .IN2(g345), .Q(n1319) );
  NOR2X1 U1549 ( .IN1(n1710), .IN2(n1022), .QN(n1992) );
  AND2X1 U1550 ( .IN1(n1805), .IN2(n1857), .Q(n1806) );
  OA21X1 U1551 ( .IN1(g119), .IN2(n1556), .IN3(g109), .Q(n2005) );
  NBUFFX2 U1552 ( .INP(g965), .Z(n1019) );
  INVX0 U1553 ( .INP(g109), .ZN(n1022) );
  XNOR3X1 U1554 ( .IN1(n1890), .IN2(n1911), .IN3(n1017), .Q(n1016) );
  XOR2X1 U1555 ( .IN1(n1769), .IN2(n1850), .Q(n1017) );
  AND2X1 U1556 ( .IN1(n1265), .IN2(n1267), .Q(n1029) );
  AND3X1 U1557 ( .IN1(n1150), .IN2(n1420), .IN3(n1418), .Q(n1018) );
  NOR2X0 U1558 ( .IN1(n1091), .IN2(n1090), .QN(n1020) );
  NAND2X0 U1559 ( .IN1(g109), .IN2(g10724), .QN(n1021) );
  NOR4X0 U1560 ( .IN1(n1877), .IN2(n1876), .IN3(g10724), .IN4(g10719), .QN(
        n1878) );
  AO21X1 U1561 ( .IN1(n1318), .IN2(n2021), .IN3(n1319), .Q(g11625) );
  AOI22X1 U1562 ( .IN1(n1267), .IN2(n1226), .IN3(n1266), .IN4(n1029), .QN(
        g11647) );
  AO21X1 U1563 ( .IN1(n1129), .IN2(n1115), .IN3(n1022), .Q(n1420) );
  OAI21X1 U1564 ( .IN1(n1023), .IN2(n1159), .IN3(g109), .QN(n1419) );
  INVX0 U1565 ( .INP(n1167), .ZN(n1023) );
  NAND4X0 U1566 ( .IN1(n1208), .IN2(n1204), .IN3(n1205), .IN4(n1344), .QN(
        n1354) );
  OA21X1 U1567 ( .IN1(n1083), .IN2(n1082), .IN3(g109), .Q(n1098) );
  NOR3X0 U1568 ( .IN1(n1302), .IN2(n1301), .IN3(n1300), .QN(n1307) );
  INVX0 U1569 ( .INP(g1822), .ZN(n1486) );
  NOR2X0 U1570 ( .IN1(n1311), .IN2(g1317), .QN(n1331) );
  NAND2X0 U1571 ( .IN1(g18), .IN2(g115), .QN(n1556) );
  NAND2X0 U1572 ( .IN1(n1289), .IN2(n1288), .QN(n1311) );
  INVX0 U1573 ( .INP(n1910), .ZN(n1289) );
  NAND2X0 U1574 ( .IN1(g1814), .IN2(n1486), .QN(n1592) );
  INVX0 U1575 ( .INP(n1313), .ZN(n1314) );
  NAND2X0 U1576 ( .IN1(g1336), .IN2(g11561), .QN(n1521) );
  NAND2X0 U1577 ( .IN1(n1286), .IN2(n1331), .QN(n1306) );
  NAND2X0 U1578 ( .IN1(n1331), .IN2(n1303), .QN(n1304) );
  INVX0 U1579 ( .INP(n1307), .ZN(n1303) );
  XNOR3X1 U1580 ( .IN1(n1360), .IN2(g10664), .IN3(g10722), .Q(n2026) );
  MUX21X1 U1581 ( .IN1(n1212), .IN2(g305), .S(n1261), .Q(n1313) );
  NAND2X0 U1582 ( .IN1(n1192), .IN2(g1727), .QN(n1343) );
  NAND2X0 U1583 ( .IN1(n1207), .IN2(g956), .QN(n1345) );
  NAND2X0 U1584 ( .IN1(n1206), .IN2(g1531), .QN(n1346) );
  NOR2X0 U1585 ( .IN1(n1052), .IN2(n1056), .QN(n1206) );
  NAND4X0 U1586 ( .IN1(n1940), .IN2(n1945), .IN3(n1778), .IN4(n1942), .QN(
        n1694) );
  NOR2X0 U1587 ( .IN1(g12), .IN2(n1556), .QN(n1710) );
  NAND3X0 U1588 ( .IN1(n1733), .IN2(g1840), .IN3(n1591), .QN(n1851) );
  INVX0 U1589 ( .INP(g1834), .ZN(n1591) );
  INVX0 U1590 ( .INP(g1828), .ZN(n1788) );
  INVX0 U1591 ( .INP(g605), .ZN(n1942) );
  INVX0 U1592 ( .INP(g599), .ZN(n1778) );
  MUX21X1 U1593 ( .IN1(n1251), .IN2(g333), .S(n1261), .Q(n1752) );
  INVX0 U1594 ( .INP(g591), .ZN(n1940) );
  NAND2X0 U1595 ( .IN1(n1245), .IN2(g309), .QN(n1236) );
  NOR2X0 U1596 ( .IN1(n1223), .IN2(n1092), .QN(n1187) );
  NOR2X0 U1597 ( .IN1(g1868), .IN2(n1375), .QN(n1733) );
  NAND4X0 U1598 ( .IN1(n1487), .IN2(n1591), .IN3(n1486), .IN4(n1788), .QN(
        n1903) );
  INVX0 U1599 ( .INP(g611), .ZN(n1945) );
  NAND2X0 U1600 ( .IN1(g798), .IN2(g794), .QN(n1957) );
  NAND2X0 U1601 ( .IN1(n1287), .IN2(n1636), .QN(n1910) );
  NOR2X0 U1602 ( .IN1(g1703), .IN2(n1699), .QN(n1881) );
  NAND2X0 U1603 ( .IN1(g1703), .IN2(g1696), .QN(n1913) );
  NAND2X0 U1604 ( .IN1(g48), .IN2(n1362), .QN(n2024) );
  NOR2X0 U1605 ( .IN1(n1804), .IN2(n1915), .QN(n1916) );
  NAND2X0 U1606 ( .IN1(n1590), .IN2(n1379), .QN(n1828) );
  INVX0 U1607 ( .INP(g1713), .ZN(n1636) );
  NAND2X0 U1608 ( .IN1(g1703), .IN2(n1699), .QN(n1978) );
  NOR2X0 U1609 ( .IN1(n1022), .IN2(n1289), .QN(n2010) );
  INVX0 U1610 ( .INP(n2007), .ZN(n1971) );
  INVX0 U1611 ( .INP(n1978), .ZN(n2006) );
  NOR2X0 U1612 ( .IN1(n1961), .IN2(n2004), .QN(n2003) );
  INVX0 U1613 ( .INP(n1871), .ZN(n1986) );
  NOR2X0 U1614 ( .IN1(n1961), .IN2(n1726), .QN(n1991) );
  NOR2X0 U1615 ( .IN1(n1732), .IN2(n1804), .QN(n2002) );
  MUX21X1 U1616 ( .IN1(g1448), .IN2(g1607), .S(n1992), .Q(g6515) );
  MUX21X1 U1617 ( .IN1(g956), .IN2(g845), .S(n1934), .Q(g11306) );
  AND2X1 U1618 ( .IN1(n1332), .IN2(n1312), .Q(g11561) );
  MUX21X1 U1619 ( .IN1(g1486), .IN2(g1540), .S(n1992), .Q(g6541) );
  NAND4X0 U1620 ( .IN1(n1329), .IN2(n1328), .IN3(n1325), .IN4(n1327), .QN(
        g10664) );
  MUX21X1 U1621 ( .IN1(g1814), .IN2(n1487), .S(n1493), .Q(n1494) );
  MUX21X1 U1622 ( .IN1(n1330), .IN2(g363), .S(n2008), .Q(g11486) );
  MUX21X1 U1623 ( .IN1(n1324), .IN2(g357), .S(n2008), .Q(g11484) );
  NAND2X0 U1624 ( .IN1(n1332), .IN2(n1030), .QN(n1309) );
  NAND2X0 U1625 ( .IN1(n1306), .IN2(n1305), .QN(n1310) );
  MUX21X1 U1626 ( .IN1(g1499), .IN2(g1531), .S(n1992), .Q(g6528) );
  MUX21X1 U1627 ( .IN1(g962), .IN2(g853), .S(n1934), .Q(g11310) );
  MUX21X1 U1628 ( .IN1(g1520), .IN2(g1571), .S(n1992), .Q(g6469) );
  MUX21X1 U1629 ( .IN1(g170), .IN2(g284), .S(n2005), .Q(g6934) );
  MUX21X1 U1630 ( .IN1(n1613), .IN2(n1612), .S(g981), .Q(g11392) );
  NOR2X0 U1631 ( .IN1(n1747), .IN2(n1746), .QN(n1934) );
  INVX0 U1632 ( .INP(n2009), .ZN(n1024) );
  INVX0 U1633 ( .INP(n1024), .ZN(n1025) );
  MUX21X1 U1634 ( .IN1(g330), .IN2(n1262), .S(n1211), .Q(n1330) );
  MUX21X1 U1635 ( .IN1(g315), .IN2(n1253), .S(n1453), .Q(n2009) );
  NAND4X0 U1636 ( .IN1(n1018), .IN2(n1419), .IN3(n1876), .IN4(n1209), .QN(
        n1027) );
  MUX21X1 U1637 ( .IN1(g944), .IN2(g829), .S(n1934), .Q(g11298) );
  NBUFFX2 U1638 ( .INP(n2010), .Z(n1028) );
  XNOR3X1 U1639 ( .IN1(n1769), .IN2(n1850), .IN3(n1264), .Q(n1316) );
  INVX0 U1640 ( .INP(g1814), .ZN(n1487) );
  INVX0 U1641 ( .INP(n2021), .ZN(n2008) );
  NOR2X0 U1642 ( .IN1(n2020), .IN2(g754), .QN(n2021) );
  AND2X1 U1643 ( .IN1(n1331), .IN2(g1796), .Q(n1030) );
  INVX0 U1644 ( .INP(n1276), .ZN(n1838) );
  AO22X1 U1645 ( .IN1(n1188), .IN2(g12), .IN3(n1185), .IN4(g4), .Q(n1031) );
  AND2X1 U1646 ( .IN1(g1027), .IN2(g1032), .Q(n1032) );
  INVX0 U1647 ( .INP(n1763), .ZN(n1288) );
  NOR4X0 U1648 ( .IN1(g486), .IN2(g491), .IN3(g511), .IN4(g538), .QN(n1034) );
  NOR4X0 U1649 ( .IN1(g501), .IN2(g496), .IN3(g542), .IN4(g534), .QN(n1033) );
  INVX0 U1650 ( .INP(g476), .ZN(n1238) );
  INVX0 U1651 ( .INP(g506), .ZN(n1260) );
  NAND4X0 U1652 ( .IN1(n1034), .IN2(n1033), .IN3(n1238), .IN4(n1260), .QN(
        n1035) );
  NOR4X0 U1653 ( .IN1(g516), .IN2(g481), .IN3(g530), .IN4(n1035), .QN(n1036)
         );
  NOR2X0 U1654 ( .IN1(n1036), .IN2(g521), .QN(n1037) );
  MUX21X1 U1655 ( .IN1(n1037), .IN2(g521), .S(g525), .Q(n1981) );
  INVX0 U1656 ( .INP(g456), .ZN(n1469) );
  NOR4X0 U1657 ( .IN1(g461), .IN2(g471), .IN3(g466), .IN4(n1469), .QN(n1038)
         );
  XOR2X1 U1658 ( .IN1(n1981), .IN2(n1038), .Q(n1212) );
  OR4X1 U1659 ( .IN1(g841), .IN2(g829), .IN3(g853), .IN4(g837), .Q(n1039) );
  OR4X1 U1660 ( .IN1(g849), .IN2(g857), .IN3(g833), .IN4(n1039), .Q(n1043) );
  INVX0 U1661 ( .INP(g861), .ZN(n1041) );
  INVX0 U1662 ( .INP(g845), .ZN(n1040) );
  NAND2X0 U1663 ( .IN1(n1041), .IN2(n1040), .QN(n1042) );
  NOR2X0 U1664 ( .IN1(n1043), .IN2(n1042), .QN(n1257) );
  INVX0 U1665 ( .INP(g42), .ZN(n1223) );
  INVX0 U1666 ( .INP(g31), .ZN(n1362) );
  NOR2X0 U1667 ( .IN1(g41), .IN2(n2024), .QN(n1060) );
  NOR2X0 U1668 ( .IN1(g46), .IN2(g47), .QN(n1224) );
  NAND2X0 U1669 ( .IN1(n1060), .IN2(n1224), .QN(n1095) );
  INVX0 U1670 ( .INP(n1095), .ZN(n1101) );
  INVX0 U1671 ( .INP(g43), .ZN(n1051) );
  INVX0 U1672 ( .INP(g45), .ZN(n1220) );
  NAND4X0 U1673 ( .IN1(g44), .IN2(n1101), .IN3(n1051), .IN4(n1220), .QN(n1092)
         );
  NAND2X0 U1674 ( .IN1(n1187), .IN2(g281), .QN(n1046) );
  NAND2X0 U1675 ( .IN1(g44), .IN2(g43), .QN(n1044) );
  NOR2X0 U1676 ( .IN1(g45), .IN2(n1044), .QN(n1047) );
  NAND2X0 U1677 ( .IN1(n1223), .IN2(n1047), .QN(n1100) );
  INVX0 U1678 ( .INP(n1100), .ZN(n1052) );
  NAND2X0 U1679 ( .IN1(n1047), .IN2(n1101), .QN(n1056) );
  NAND2X0 U1680 ( .IN1(n1206), .IN2(g1543), .QN(n1045) );
  NAND2X0 U1681 ( .IN1(n1046), .IN2(n1045), .QN(n1067) );
  NAND2X0 U1682 ( .IN1(g39), .IN2(n2024), .QN(n1065) );
  INVX0 U1683 ( .INP(g47), .ZN(n1059) );
  AND2X1 U1684 ( .IN1(n1059), .IN2(g46), .Q(n1338) );
  NAND2X0 U1685 ( .IN1(n1060), .IN2(n1338), .QN(n1072) );
  INVX0 U1686 ( .INP(n1072), .ZN(n1053) );
  NOR2X0 U1687 ( .IN1(g44), .IN2(n1051), .QN(n1102) );
  NAND4X0 U1688 ( .IN1(n1053), .IN2(g42), .IN3(g45), .IN4(n1102), .QN(n1118)
         );
  NAND4X0 U1689 ( .IN1(n1053), .IN2(g42), .IN3(g45), .IN4(n1051), .QN(n1048)
         );
  NAND4X0 U1690 ( .IN1(n1060), .IN2(g46), .IN3(g47), .IN4(n1052), .QN(n1107)
         );
  NAND2X0 U1691 ( .IN1(g42), .IN2(n1047), .QN(n1061) );
  NOR2X0 U1692 ( .IN1(n1072), .IN2(n1061), .QN(n1215) );
  INVX0 U1693 ( .INP(n1215), .ZN(n1121) );
  NAND4X0 U1694 ( .IN1(n1118), .IN2(n1048), .IN3(n1107), .IN4(n1121), .QN(
        n1050) );
  INVX0 U1695 ( .INP(n1092), .ZN(n1049) );
  NOR3X0 U1696 ( .IN1(n1050), .IN2(n1049), .IN3(n2024), .QN(n1054) );
  INVX0 U1697 ( .INP(g44), .ZN(n1221) );
  NAND3X0 U1698 ( .IN1(n1221), .IN2(n1051), .IN3(g45), .QN(n1055) );
  NOR2X0 U1699 ( .IN1(g42), .IN2(n1055), .QN(n1070) );
  NAND2X0 U1700 ( .IN1(n1053), .IN2(n1070), .QN(n1071) );
  NAND2X0 U1701 ( .IN1(n1053), .IN2(n1052), .QN(n1104) );
  NAND3X0 U1702 ( .IN1(n1054), .IN2(n1071), .IN3(n1104), .QN(n1058) );
  INVX0 U1703 ( .INP(n1055), .ZN(n1068) );
  NAND2X0 U1704 ( .IN1(n1068), .IN2(n1101), .QN(n1096) );
  NAND2X0 U1705 ( .IN1(n1056), .IN2(n1096), .QN(n1057) );
  NOR2X0 U1706 ( .IN1(n1058), .IN2(n1057), .QN(n1087) );
  NOR2X0 U1707 ( .IN1(g46), .IN2(n1059), .QN(n1334) );
  NAND2X0 U1708 ( .IN1(n1060), .IN2(n1334), .QN(n1099) );
  INVX0 U1709 ( .INP(n1099), .ZN(n1069) );
  NAND4X0 U1710 ( .IN1(g44), .IN2(g45), .IN3(g43), .IN4(n1069), .QN(n1086) );
  NOR2X0 U1711 ( .IN1(n1061), .IN2(n1099), .QN(n1199) );
  INVX0 U1712 ( .INP(n1199), .ZN(n1085) );
  NAND2X0 U1713 ( .IN1(n1068), .IN2(n1069), .QN(n1062) );
  NAND4X0 U1714 ( .IN1(n1087), .IN2(n1086), .IN3(n1085), .IN4(n1062), .QN(
        n1103) );
  NAND2X0 U1715 ( .IN1(n1199), .IN2(g1188), .QN(n1063) );
  AND3X1 U1716 ( .IN1(n1103), .IN2(n1107), .IN3(n1063), .Q(n1064) );
  NAND2X0 U1717 ( .IN1(n1065), .IN2(n1064), .QN(n1066) );
  NOR2X0 U1718 ( .IN1(n1067), .IN2(n1066), .QN(n1213) );
  NAND2X0 U1719 ( .IN1(g42), .IN2(n1068), .QN(n1079) );
  NOR2X0 U1720 ( .IN1(n1079), .IN2(n1099), .QN(n1196) );
  NAND2X0 U1721 ( .IN1(n1070), .IN2(n1069), .QN(n1084) );
  INVX0 U1722 ( .INP(n1084), .ZN(n1195) );
  AO22X1 U1723 ( .IN1(n1196), .IN2(g1308), .IN3(g1333), .IN4(n1195), .Q(n1074)
         );
  NOR2X0 U1724 ( .IN1(n1072), .IN2(n1079), .QN(n1183) );
  AO22X1 U1725 ( .IN1(n1207), .IN2(g968), .IN3(g944), .IN4(n1183), .Q(n1073)
         );
  NOR2X0 U1726 ( .IN1(n1074), .IN2(n1073), .QN(n1218) );
  AOI22X1 U1727 ( .IN1(n1215), .IN2(g919), .IN3(n1196), .IN4(g1311), .QN(n1329) );
  NAND3X0 U1728 ( .IN1(n1213), .IN2(n1218), .IN3(n1329), .QN(n1083) );
  NOR2X0 U1729 ( .IN1(n1223), .IN2(n1086), .QN(n1192) );
  INVX0 U1730 ( .INP(n1192), .ZN(n1075) );
  INVX0 U1731 ( .INP(n1196), .ZN(n1160) );
  NAND4X0 U1732 ( .IN1(n1087), .IN2(n1075), .IN3(n1085), .IN4(n1160), .QN(
        n1077) );
  NAND2X0 U1733 ( .IN1(n1187), .IN2(g284), .QN(n1076) );
  NAND2X0 U1734 ( .IN1(n1077), .IN2(n1076), .QN(n1078) );
  NOR2X0 U1735 ( .IN1(n1078), .IN2(n1015), .QN(n1325) );
  NOR2X0 U1736 ( .IN1(n1079), .IN2(n1095), .QN(n1214) );
  AO22X1 U1737 ( .IN1(n1215), .IN2(g916), .IN3(n1214), .IN4(g1586), .Q(n1080)
         );
  AO22X1 U1738 ( .IN1(g1191), .IN2(n1199), .IN3(g40), .IN4(n2024), .Q(n1326)
         );
  NOR2X0 U1739 ( .IN1(n1080), .IN2(n1326), .QN(n1081) );
  AOI22X1 U1740 ( .IN1(n1183), .IN2(g947), .IN3(n1214), .IN4(g1589), .QN(n1328) );
  NAND3X0 U1741 ( .IN1(n1325), .IN2(n1081), .IN3(n1328), .QN(n1082) );
  NAND2X0 U1742 ( .IN1(g278), .IN2(n1187), .QN(n1089) );
  NAND2X0 U1743 ( .IN1(n1207), .IN2(g965), .QN(n1088) );
  NAND4X0 U1744 ( .IN1(n1087), .IN2(n1086), .IN3(n1085), .IN4(n1084), .QN(
        n1136) );
  NAND3X0 U1745 ( .IN1(n1089), .IN2(n1088), .IN3(n1136), .QN(n1091) );
  AO22X1 U1746 ( .IN1(g1185), .IN2(n1199), .IN3(g38), .IN4(n2024), .Q(n1090)
         );
  NOR2X0 U1747 ( .IN1(n1091), .IN2(n1090), .QN(n1323) );
  NAND2X0 U1748 ( .IN1(n1206), .IN2(g1540), .QN(n1094) );
  NOR2X0 U1749 ( .IN1(g42), .IN2(n1092), .QN(n1186) );
  AOI22X1 U1750 ( .IN1(n1215), .IN2(g913), .IN3(n1186), .IN4(g302), .QN(n1093)
         );
  AND2X1 U1751 ( .IN1(n1094), .IN2(n1093), .Q(n1322) );
  NOR2X0 U1752 ( .IN1(n1100), .IN2(n1095), .QN(n1197) );
  AOI22X1 U1753 ( .IN1(n1214), .IN2(g1583), .IN3(n1197), .IN4(g1564), .QN(
        n1321) );
  NOR2X0 U1754 ( .IN1(g42), .IN2(n1096), .QN(n1184) );
  AOI22X1 U1755 ( .IN1(n1195), .IN2(g1330), .IN3(n1184), .IN4(g1607), .QN(
        n1320) );
  NAND4X0 U1756 ( .IN1(n1323), .IN2(n1322), .IN3(n1321), .IN4(n1320), .QN(
        n1097) );
  AND2X1 U1757 ( .IN1(n1097), .IN2(g109), .Q(n1653) );
  NOR2X0 U1758 ( .IN1(n1653), .IN2(n1098), .QN(n1150) );
  NAND2X0 U1759 ( .IN1(g950), .IN2(n1207), .QN(n1110) );
  NAND2X0 U1760 ( .IN1(n1186), .IN2(g287), .QN(n1109) );
  NOR2X0 U1761 ( .IN1(n1100), .IN2(n1099), .QN(n1198) );
  NAND3X0 U1762 ( .IN1(n1102), .IN2(n1101), .IN3(n1220), .QN(n1111) );
  INVX0 U1763 ( .INP(n1111), .ZN(n1137) );
  OR3X1 U1764 ( .IN1(n1198), .IN2(n1137), .IN3(n1103), .Q(n1193) );
  AOI22X1 U1765 ( .IN1(n1199), .IN2(g1170), .IN3(n1198), .IN4(g1194), .QN(
        n1106) );
  INVX0 U1766 ( .INP(n1104), .ZN(n1151) );
  NAND2X0 U1767 ( .IN1(n1151), .IN2(g922), .QN(n1105) );
  AND4X1 U1768 ( .IN1(n1107), .IN2(n1193), .IN3(n1106), .IN4(n1105), .Q(n1108)
         );
  AND3X1 U1769 ( .IN1(n1110), .IN2(n1109), .IN3(n1108), .Q(n1114) );
  NOR2X0 U1770 ( .IN1(g42), .IN2(n1111), .QN(n1188) );
  NOR2X0 U1771 ( .IN1(n1223), .IN2(n1111), .QN(n1185) );
  AOI22X1 U1772 ( .IN1(n1188), .IN2(g119), .IN3(n1185), .IN4(g123), .QN(n1113)
         );
  AOI22X1 U1773 ( .IN1(n1196), .IN2(g1336), .IN3(n1214), .IN4(g1567), .QN(
        n1112) );
  NAND2X0 U1774 ( .IN1(g263), .IN2(n1187), .QN(n1117) );
  NAND2X0 U1775 ( .IN1(g1549), .IN2(n1197), .QN(n1116) );
  NAND2X0 U1776 ( .IN1(n1117), .IN2(n1116), .QN(n1128) );
  NAND2X0 U1777 ( .IN1(g971), .IN2(n1183), .QN(n1124) );
  INVX0 U1778 ( .INP(g898), .ZN(n1120) );
  INVX0 U1779 ( .INP(n1118), .ZN(n1194) );
  NAND2X0 U1780 ( .IN1(g886), .IN2(n1194), .QN(n1119) );
  OA21X1 U1781 ( .IN1(n1121), .IN2(n1120), .IN3(n1119), .Q(n1123) );
  NAND2X0 U1782 ( .IN1(g1314), .IN2(n1195), .QN(n1122) );
  NAND3X0 U1783 ( .IN1(n1124), .IN2(n1123), .IN3(n1122), .QN(n1127) );
  AO22X1 U1784 ( .IN1(g1721), .IN2(n1192), .IN3(g33), .IN4(n2024), .Q(n1126)
         );
  AO22X1 U1785 ( .IN1(n1206), .IN2(g1524), .IN3(n1184), .IN4(g1592), .Q(n1125)
         );
  NOR4X0 U1786 ( .IN1(n1128), .IN2(n1127), .IN3(n1126), .IN4(n1125), .QN(n1129) );
  AOI22X1 U1787 ( .IN1(g1182), .IN2(n1199), .IN3(g37), .IN4(n2024), .QN(n1133)
         );
  NAND2X0 U1788 ( .IN1(g1327), .IN2(n1195), .QN(n1131) );
  NAND2X0 U1789 ( .IN1(g910), .IN2(n1215), .QN(n1130) );
  AND2X1 U1790 ( .IN1(n1131), .IN2(n1130), .Q(n1132) );
  NAND2X0 U1791 ( .IN1(n1133), .IN2(n1132), .QN(n1134) );
  INVX0 U1792 ( .INP(n1134), .ZN(n1149) );
  AO22X1 U1793 ( .IN1(n1187), .IN2(g275), .IN3(n1214), .IN4(g1580), .Q(n1135)
         );
  AOI21X1 U1794 ( .IN1(n1207), .IN2(g962), .IN3(n1135), .QN(n1148) );
  NAND2X0 U1795 ( .IN1(g1561), .IN2(n1197), .QN(n1141) );
  NAND2X0 U1796 ( .IN1(g7), .IN2(n1185), .QN(n1140) );
  NAND2X0 U1797 ( .IN1(g16), .IN2(n1188), .QN(n1139) );
  OR2X1 U1798 ( .IN1(n1137), .IN2(n1136), .Q(n1138) );
  NAND4X0 U1799 ( .IN1(n1141), .IN2(n1140), .IN3(n1139), .IN4(n1138), .QN(
        n1143) );
  AND2X1 U1800 ( .IN1(g1604), .IN2(n1184), .Q(n1142) );
  NOR2X0 U1801 ( .IN1(n1143), .IN2(n1142), .QN(n1147) );
  AND2X1 U1802 ( .IN1(n1186), .IN2(g299), .Q(n1145) );
  AO22X1 U1803 ( .IN1(n1192), .IN2(g1733), .IN3(n1206), .IN4(g1537), .Q(n1144)
         );
  NOR2X0 U1804 ( .IN1(n1145), .IN2(n1144), .QN(n1146) );
  NAND4X0 U1805 ( .IN1(n1149), .IN2(n1147), .IN3(n1148), .IN4(n1146), .QN(
        g10724) );
  NAND2X0 U1806 ( .IN1(g109), .IN2(g10724), .QN(n1418) );
  AND3X1 U1807 ( .IN1(n1150), .IN2(n1420), .IN3(n1418), .Q(n1210) );
  AOI22X1 U1808 ( .IN1(g1571), .IN2(n1214), .IN3(g34), .IN4(n2024), .QN(n1158)
         );
  AO22X1 U1809 ( .IN1(n1206), .IN2(g1528), .IN3(n1184), .IN4(g1595), .Q(n1155)
         );
  AO22X1 U1810 ( .IN1(n1207), .IN2(g953), .IN3(n1197), .IN4(g1552), .Q(n1154)
         );
  AO22X1 U1811 ( .IN1(n1151), .IN2(g925), .IN3(n1194), .IN4(g889), .Q(n1153)
         );
  AND2X1 U1812 ( .IN1(g1318), .IN2(n1195), .Q(n1152) );
  NOR4X0 U1813 ( .IN1(n1155), .IN2(n1154), .IN3(n1153), .IN4(n1152), .QN(n1157) );
  NAND2X0 U1814 ( .IN1(n1192), .IN2(g1724), .QN(n1156) );
  NAND4X0 U1815 ( .IN1(n1158), .IN2(n1157), .IN3(n1193), .IN4(n1156), .QN(
        n1159) );
  INVX0 U1816 ( .INP(n1159), .ZN(n1168) );
  INVX0 U1817 ( .INP(g1341), .ZN(n1507) );
  NOR2X0 U1818 ( .IN1(n1160), .IN2(n1507), .QN(n1166) );
  NAND2X0 U1819 ( .IN1(n1183), .IN2(g976), .QN(n1163) );
  NAND2X0 U1820 ( .IN1(n1186), .IN2(g290), .QN(n1162) );
  AOI22X1 U1821 ( .IN1(n1199), .IN2(g1173), .IN3(n1198), .IN4(g1197), .QN(
        n1161) );
  NAND3X0 U1822 ( .IN1(n1163), .IN2(n1162), .IN3(n1161), .QN(n1165) );
  AO22X1 U1823 ( .IN1(n1215), .IN2(g901), .IN3(n1187), .IN4(g266), .Q(n1164)
         );
  NOR4X0 U1824 ( .IN1(n1166), .IN2(n1165), .IN3(n1164), .IN4(n1031), .QN(n1167) );
  NAND2X0 U1825 ( .IN1(n1168), .IN2(n1167), .QN(g10720) );
  AO22X1 U1826 ( .IN1(n1215), .IN2(g907), .IN3(n1214), .IN4(g1577), .Q(n1172)
         );
  AO22X1 U1827 ( .IN1(n1194), .IN2(g895), .IN3(n1197), .IN4(g1558), .Q(n1171)
         );
  AO22X1 U1828 ( .IN1(n1199), .IN2(g1179), .IN3(n1198), .IN4(g1203), .Q(n1170)
         );
  AO22X1 U1829 ( .IN1(n1196), .IN2(g1351), .IN3(n1195), .IN4(g1324), .Q(n1169)
         );
  NOR4X0 U1830 ( .IN1(n1172), .IN2(n1171), .IN3(n1170), .IN4(n1169), .QN(n1182) );
  NAND2X0 U1831 ( .IN1(n1187), .IN2(g272), .QN(n1181) );
  AO22X1 U1832 ( .IN1(n1206), .IN2(g1534), .IN3(n1184), .IN4(g1601), .Q(n1175)
         );
  AO22X1 U1833 ( .IN1(g959), .IN2(n1207), .IN3(g36), .IN4(n2024), .Q(n1174) );
  AO22X1 U1834 ( .IN1(n1188), .IN2(g17), .IN3(n1185), .IN4(g8), .Q(n1173) );
  NOR3X0 U1835 ( .IN1(n1175), .IN2(n1174), .IN3(n1173), .QN(n1180) );
  NAND2X0 U1836 ( .IN1(g986), .IN2(n1183), .QN(n1178) );
  NAND2X0 U1837 ( .IN1(g1730), .IN2(n1192), .QN(n1177) );
  NAND2X0 U1838 ( .IN1(n1186), .IN2(g296), .QN(n1176) );
  NAND4X0 U1839 ( .IN1(n1182), .IN2(n1181), .IN3(n1180), .IN4(n1179), .QN(
        g10722) );
  AOI22X1 U1840 ( .IN1(g981), .IN2(n1183), .IN3(g35), .IN4(n2024), .QN(n1349)
         );
  AOI22X1 U1841 ( .IN1(n1185), .IN2(g1), .IN3(n1184), .IN4(g1598), .QN(n1348)
         );
  NAND2X0 U1842 ( .IN1(n1186), .IN2(g293), .QN(n1191) );
  NAND2X0 U1843 ( .IN1(n1187), .IN2(g269), .QN(n1190) );
  NAND2X0 U1844 ( .IN1(n1188), .IN2(g9), .QN(n1189) );
  AND3X1 U1845 ( .IN1(n1191), .IN2(n1190), .IN3(n1189), .Q(n1347) );
  AND3X1 U1846 ( .IN1(n1349), .IN2(n1348), .IN3(n1347), .Q(n1205) );
  AND2X1 U1847 ( .IN1(n1343), .IN2(n1193), .Q(n1204) );
  AO22X1 U1848 ( .IN1(n1194), .IN2(g892), .IN3(n1214), .IN4(g1574), .Q(n1203)
         );
  AO22X1 U1849 ( .IN1(n1196), .IN2(g1346), .IN3(n1195), .IN4(g1321), .Q(n1202)
         );
  AO22X1 U1850 ( .IN1(n1215), .IN2(g904), .IN3(n1197), .IN4(g1555), .Q(n1201)
         );
  AO22X1 U1851 ( .IN1(n1199), .IN2(g1176), .IN3(n1198), .IN4(g1200), .Q(n1200)
         );
  NOR4X0 U1852 ( .IN1(n1203), .IN2(n1202), .IN3(n1201), .IN4(n1200), .QN(n1344) );
  AND2X1 U1853 ( .IN1(n1346), .IN2(n1345), .Q(n1208) );
  AND2X1 U1854 ( .IN1(n1354), .IN2(g109), .Q(n1333) );
  INVX0 U1855 ( .INP(n1333), .ZN(n1209) );
  NAND4X0 U1856 ( .IN1(n1210), .IN2(n1419), .IN3(n1876), .IN4(n1209), .QN(
        n1256) );
  NAND2X0 U1857 ( .IN1(n1257), .IN2(n1256), .QN(n1211) );
  INVX0 U1858 ( .INP(n1250), .ZN(n1245) );
  INVX0 U1859 ( .INP(n1026), .ZN(n1467) );
  INVX0 U1860 ( .INP(n1213), .ZN(n1217) );
  AO22X1 U1861 ( .IN1(n1215), .IN2(g916), .IN3(n1214), .IN4(g1586), .Q(n1216)
         );
  NOR2X0 U1862 ( .IN1(n1217), .IN2(n1216), .QN(n1219) );
  NAND2X0 U1863 ( .IN1(n1219), .IN2(n1218), .QN(g10663) );
  NOR4X0 U1864 ( .IN1(g48), .IN2(g41), .IN3(g43), .IN4(g30), .QN(n1222) );
  NAND3X0 U1865 ( .IN1(n1222), .IN2(n1221), .IN3(n1220), .QN(n1336) );
  NOR2X0 U1866 ( .IN1(n1223), .IN2(n1336), .QN(n1335) );
  AND2X1 U1867 ( .IN1(n1224), .IN2(n1335), .Q(n1877) );
  OR2X1 U1868 ( .IN1(g10663), .IN2(n1877), .Q(n1276) );
  NAND2X0 U1869 ( .IN1(n1313), .IN2(n1838), .QN(n1265) );
  NAND2X0 U1870 ( .IN1(n1265), .IN2(n1838), .QN(n1225) );
  INVX0 U1871 ( .INP(g750), .ZN(n2020) );
  NAND2X0 U1872 ( .IN1(n1225), .IN2(n2021), .QN(n1226) );
  NAND2X0 U1873 ( .IN1(n1026), .IN2(g327), .QN(n1231) );
  INVX0 U1874 ( .INP(g501), .ZN(n1228) );
  INVX0 U1875 ( .INP(g471), .ZN(n1468) );
  NAND4X0 U1876 ( .IN1(g461), .IN2(g466), .IN3(n1468), .IN4(n1469), .QN(n1227)
         );
  MUX21X1 U1877 ( .IN1(n1228), .IN2(g501), .S(n1227), .Q(n1229) );
  NAND2X0 U1878 ( .IN1(n1229), .IN2(n1467), .QN(n1230) );
  NAND2X0 U1879 ( .IN1(n1231), .IN2(n1230), .QN(n1911) );
  INVX0 U1880 ( .INP(g516), .ZN(n1233) );
  INVX0 U1881 ( .INP(g461), .ZN(n1512) );
  INVX0 U1882 ( .INP(g466), .ZN(n1730) );
  NAND4X0 U1883 ( .IN1(g456), .IN2(g471), .IN3(n1512), .IN4(n1730), .QN(n1232)
         );
  MUX21X1 U1884 ( .IN1(n1233), .IN2(g516), .S(n1232), .Q(n1234) );
  NAND2X0 U1885 ( .IN1(n1467), .IN2(n1234), .QN(n1235) );
  NAND2X0 U1886 ( .IN1(n1236), .IN2(n1235), .QN(n1890) );
  NAND4X0 U1887 ( .IN1(g461), .IN2(g471), .IN3(n1469), .IN4(n1730), .QN(n1237)
         );
  MUX21X1 U1888 ( .IN1(n1238), .IN2(g476), .S(n1237), .Q(n1239) );
  INVX0 U1889 ( .INP(g486), .ZN(n1241) );
  NAND4X0 U1890 ( .IN1(g456), .IN2(g461), .IN3(n1468), .IN4(n1730), .QN(n1240)
         );
  MUX21X1 U1891 ( .IN1(n1241), .IN2(g486), .S(n1240), .Q(n1242) );
  MUX21X1 U1892 ( .IN1(n1242), .IN2(g318), .S(n1245), .Q(n1850) );
  INVX0 U1893 ( .INP(g491), .ZN(n1244) );
  NOR4X0 U1894 ( .IN1(g461), .IN2(g456), .IN3(g471), .IN4(n1730), .QN(n1243)
         );
  MUX21X1 U1895 ( .IN1(g491), .IN2(n1244), .S(n1243), .Q(n1246) );
  MUX21X1 U1896 ( .IN1(n1246), .IN2(g321), .S(n1245), .Q(n1830) );
  INVX0 U1897 ( .INP(g511), .ZN(n1249) );
  NAND3X0 U1898 ( .IN1(g471), .IN2(n1512), .IN3(n1730), .QN(n1247) );
  NOR2X0 U1899 ( .IN1(g456), .IN2(n1247), .QN(n1248) );
  MUX21X1 U1900 ( .IN1(g511), .IN2(n1249), .S(n1248), .Q(n1251) );
  NAND2X0 U1901 ( .IN1(n1257), .IN2(n1256), .QN(n1250) );
  INVX0 U1902 ( .INP(n1211), .ZN(n1261) );
  INVX0 U1903 ( .INP(g481), .ZN(n1980) );
  NOR4X0 U1904 ( .IN1(g471), .IN2(g456), .IN3(g466), .IN4(n1512), .QN(n1252)
         );
  MUX21X1 U1905 ( .IN1(g481), .IN2(n1980), .S(n1252), .Q(n1253) );
  NAND2X0 U1906 ( .IN1(n1257), .IN2(n1027), .QN(n1453) );
  INVX0 U1907 ( .INP(g496), .ZN(n1255) );
  NAND4X0 U1908 ( .IN1(g456), .IN2(g466), .IN3(n1512), .IN4(n1468), .QN(n1254)
         );
  MUX21X1 U1909 ( .IN1(n1255), .IN2(g496), .S(n1254), .Q(n1258) );
  NAND2X0 U1910 ( .IN1(n1257), .IN2(n1027), .QN(n1415) );
  MUX21X1 U1911 ( .IN1(g324), .IN2(n1258), .S(n1415), .Q(n1324) );
  NAND3X0 U1912 ( .IN1(g461), .IN2(g456), .IN3(g466), .QN(n1562) );
  NOR2X0 U1913 ( .IN1(g471), .IN2(n1562), .QN(n1259) );
  MUX21X1 U1914 ( .IN1(g506), .IN2(n1260), .S(n1259), .Q(n1262) );
  XNOR3X1 U1915 ( .IN1(n2009), .IN2(n1324), .IN3(n1330), .Q(n1263) );
  XNOR3X1 U1916 ( .IN1(n1830), .IN2(n1752), .IN3(n1263), .Q(n1264) );
  NAND2X0 U1917 ( .IN1(n2008), .IN2(g336), .QN(n1267) );
  NOR2X0 U1918 ( .IN1(g1280), .IN2(g1284), .QN(n1272) );
  INVX0 U1919 ( .INP(g1265), .ZN(n1292) );
  INVX0 U1920 ( .INP(g1260), .ZN(n1299) );
  INVX0 U1921 ( .INP(g1240), .ZN(n1279) );
  INVX0 U1922 ( .INP(g1270), .ZN(n1280) );
  NAND4X0 U1923 ( .IN1(n1292), .IN2(n1299), .IN3(n1279), .IN4(n1280), .QN(
        n1270) );
  OR4X1 U1924 ( .IN1(g1255), .IN2(g1250), .IN3(g1245), .IN4(g1296), .Q(n1268)
         );
  OR4X1 U1925 ( .IN1(g1235), .IN2(g1275), .IN3(g1304), .IN4(n1268), .Q(n1269)
         );
  OR4X1 U1926 ( .IN1(g1300), .IN2(g1292), .IN3(n1270), .IN4(n1269), .Q(n1271)
         );
  NAND4X0 U1927 ( .IN1(g1227), .IN2(g1223), .IN3(g1218), .IN4(g1231), .QN(
        n1763) );
  AO221X1 U1928 ( .IN1(g1284), .IN2(g1280), .IN3(n1272), .IN4(n1271), .IN5(
        n1763), .Q(n1764) );
  NAND2X0 U1929 ( .IN1(g10663), .IN2(g1032), .QN(n1275) );
  INVX0 U1930 ( .INP(g1027), .ZN(n1832) );
  NAND2X0 U1931 ( .IN1(g1032), .IN2(n1877), .QN(n1273) );
  NAND2X0 U1932 ( .IN1(n1275), .IN2(n1274), .QN(n1278) );
  NAND2X0 U1933 ( .IN1(n1276), .IN2(n1032), .QN(n1277) );
  NAND2X0 U1934 ( .IN1(n1278), .IN2(n1277), .QN(n1765) );
  XNOR2X1 U1935 ( .IN1(n1764), .IN2(n1765), .Q(n1285) );
  MUX21X1 U1936 ( .IN1(n1279), .IN2(g1240), .S(g1003), .Q(n1284) );
  MUX21X1 U1937 ( .IN1(n1280), .IN2(g1270), .S(g1023), .Q(n1283) );
  INVX0 U1938 ( .INP(g1245), .ZN(n1281) );
  MUX21X1 U1939 ( .IN1(n1281), .IN2(g1245), .S(g999), .Q(n1282) );
  NAND4X0 U1940 ( .IN1(n1285), .IN2(n1284), .IN3(n1283), .IN4(n1282), .QN(
        n1286) );
  INVX0 U1941 ( .INP(n1286), .ZN(n1308) );
  NOR2X0 U1942 ( .IN1(g1703), .IN2(g1696), .QN(n1287) );
  INVX0 U1943 ( .INP(g1235), .ZN(n1290) );
  MUX21X1 U1944 ( .IN1(n1290), .IN2(g1235), .S(g991), .Q(n1297) );
  INVX0 U1945 ( .INP(g1275), .ZN(n1291) );
  MUX21X1 U1946 ( .IN1(n1291), .IN2(g1275), .S(g995), .Q(n1296) );
  MUX21X1 U1947 ( .IN1(n1292), .IN2(g1265), .S(g1015), .Q(n1295) );
  INVX0 U1948 ( .INP(g1255), .ZN(n1293) );
  MUX21X1 U1949 ( .IN1(n1293), .IN2(g1255), .S(g1007), .Q(n1294) );
  NAND4X0 U1950 ( .IN1(n1297), .IN2(n1296), .IN3(n1295), .IN4(n1294), .QN(
        n1302) );
  INVX0 U1951 ( .INP(g1250), .ZN(n1298) );
  MUX21X1 U1952 ( .IN1(g1250), .IN2(n1298), .S(g1011), .Q(n1301) );
  MUX21X1 U1953 ( .IN1(g1260), .IN2(n1299), .S(g1019), .Q(n1300) );
  NAND2X0 U1954 ( .IN1(n1308), .IN2(n1307), .QN(n1332) );
  NAND2X0 U1955 ( .IN1(n1310), .IN2(n1309), .QN(g11608) );
  INVX0 U1956 ( .INP(n1311), .ZN(n1312) );
  XOR2X1 U1957 ( .IN1(n1911), .IN2(n1890), .Q(n1315) );
  XOR2X1 U1958 ( .IN1(n1315), .IN2(n1314), .Q(n1317) );
  XOR2X1 U1959 ( .IN1(n1317), .IN2(n1316), .Q(n1318) );
  NAND4X0 U1960 ( .IN1(n1020), .IN2(n1322), .IN3(n1321), .IN4(n1320), .QN(
        n2029) );
  INVX0 U1961 ( .INP(n1326), .ZN(n1327) );
  MUX21X1 U1962 ( .IN1(g1490), .IN2(g1537), .S(n1992), .Q(g6537) );
  NAND2X0 U1963 ( .IN1(n1332), .IN2(n1331), .QN(n1965) );
  MUX21X1 U1964 ( .IN1(g1776), .IN2(g1314), .S(n1965), .Q(g11604) );
  MUX21X1 U1965 ( .IN1(n1333), .IN2(g1727), .S(n1913), .Q(g10773) );
  NAND2X0 U1966 ( .IN1(n1334), .IN2(n1335), .QN(n1010) );
  NAND2X0 U1967 ( .IN1(n1338), .IN2(n1335), .QN(n1013) );
  NOR2X0 U1968 ( .IN1(g42), .IN2(n1336), .QN(n1337) );
  NAND2X0 U1969 ( .IN1(n1338), .IN2(n1337), .QN(n1012) );
  INVX0 U1970 ( .INP(g10719), .ZN(n1339) );
  NOR2X0 U1971 ( .IN1(g30), .IN2(n2024), .QN(n1361) );
  NAND2X0 U1972 ( .IN1(n1339), .IN2(n1361), .QN(g10402) );
  INVX0 U1973 ( .INP(g10664), .ZN(n1340) );
  NAND2X0 U1974 ( .IN1(n1340), .IN2(n1361), .QN(g10339) );
  INVX0 U1975 ( .INP(g10663), .ZN(n1352) );
  NAND2X0 U1976 ( .IN1(n1352), .IN2(n1361), .QN(g10336) );
  INVX0 U1977 ( .INP(g10722), .ZN(n1341) );
  NAND2X0 U1978 ( .IN1(n1341), .IN2(n1361), .QN(g10411) );
  INVX0 U1979 ( .INP(g10724), .ZN(n1342) );
  NAND2X0 U1980 ( .IN1(n1342), .IN2(n1361), .QN(g10414) );
  INVX0 U1981 ( .INP(n2029), .ZN(n1359) );
  NAND2X0 U1982 ( .IN1(n1359), .IN2(n1361), .QN(g10417) );
  INVX0 U1983 ( .INP(g10720), .ZN(n1880) );
  NAND2X0 U1984 ( .IN1(n1880), .IN2(n1361), .QN(g10405) );
  NOR2X0 U1985 ( .IN1(n1351), .IN2(n1350), .QN(n1353) );
  NAND2X0 U1986 ( .IN1(n1353), .IN2(n1352), .QN(n1356) );
  NAND2X0 U1987 ( .IN1(g10663), .IN2(n1354), .QN(n1355) );
  NAND2X0 U1988 ( .IN1(n1356), .IN2(n1355), .QN(n1357) );
  XNOR3X1 U1989 ( .IN1(n1357), .IN2(g10719), .IN3(g10720), .Q(n1358) );
  XOR3X1 U1990 ( .IN1(n1359), .IN2(g10724), .IN3(n1358), .Q(n1360) );
  NAND2X0 U1991 ( .IN1(n1361), .IN2(n2026), .QN(g10712) );
  INVX0 U1992 ( .INP(n1354), .ZN(n1879) );
  NAND2X0 U1993 ( .IN1(n1879), .IN2(n1361), .QN(g10408) );
  NOR2X0 U1994 ( .IN1(g41), .IN2(g30), .QN(n1363) );
  NAND2X0 U1995 ( .IN1(n1363), .IN2(n1362), .QN(g9931) );
  NAND3X0 U1996 ( .IN1(g109), .IN2(g746), .IN3(g745), .QN(n1817) );
  INVX0 U1997 ( .INP(n1817), .ZN(n1675) );
  NAND2X0 U1998 ( .IN1(g794), .IN2(n1675), .QN(g5849) );
  INVX0 U1999 ( .INP(g1845), .ZN(n1717) );
  NOR2X0 U2000 ( .IN1(g1822), .IN2(g1828), .QN(n1892) );
  OA21X1 U2001 ( .IN1(g1834), .IN2(n1892), .IN3(n1487), .Q(n1007) );
  INVX0 U2002 ( .INP(n1007), .ZN(n1727) );
  NAND2X0 U2003 ( .IN1(n1717), .IN2(n1727), .QN(g6755) );
  NAND2X0 U2004 ( .IN1(g18), .IN2(g225), .QN(n1666) );
  OA21X1 U2005 ( .IN1(g18), .IN2(g1624), .IN3(n1666), .Q(n1692) );
  INVX0 U2006 ( .INP(n1692), .ZN(n1690) );
  NAND2X0 U2007 ( .IN1(n1690), .IN2(n2007), .QN(n1364) );
  NOR2X0 U2008 ( .IN1(g1718), .IN2(n1364), .QN(n1783) );
  INVX0 U2009 ( .INP(n1783), .ZN(n1366) );
  NAND2X0 U2010 ( .IN1(n1971), .IN2(g1684), .QN(n1365) );
  NAND2X0 U2011 ( .IN1(n1366), .IN2(n1365), .QN(g10866) );
  INVX0 U2012 ( .INP(g1618), .ZN(n1367) );
  NAND2X0 U2013 ( .IN1(g18), .IN2(g186), .QN(n1495) );
  OA21X1 U2014 ( .IN1(g18), .IN2(n1367), .IN3(n1495), .Q(n1661) );
  INVX0 U2015 ( .INP(n1661), .ZN(n1659) );
  NAND2X0 U2016 ( .IN1(n1659), .IN2(n2007), .QN(n1368) );
  NOR2X0 U2017 ( .IN1(g1718), .IN2(n1368), .QN(n1843) );
  INVX0 U2018 ( .INP(n1843), .ZN(n1370) );
  NAND2X0 U2019 ( .IN1(n1971), .IN2(g546), .QN(n1369) );
  NAND2X0 U2020 ( .IN1(n1370), .IN2(n1369), .QN(g10791) );
  INVX0 U2021 ( .INP(g1621), .ZN(n1371) );
  NAND2X0 U2022 ( .IN1(g18), .IN2(g219), .QN(n1696) );
  OA21X1 U2023 ( .IN1(g18), .IN2(n1371), .IN3(n1696), .Q(n1537) );
  INVX0 U2024 ( .INP(n1537), .ZN(n1535) );
  NAND2X0 U2025 ( .IN1(n1535), .IN2(n2007), .QN(n1372) );
  NOR2X0 U2026 ( .IN1(g1718), .IN2(n1372), .QN(n1748) );
  INVX0 U2027 ( .INP(n1748), .ZN(n1374) );
  NAND2X0 U2028 ( .IN1(n1971), .IN2(g560), .QN(n1373) );
  NAND2X0 U2029 ( .IN1(n1374), .IN2(n1373), .QN(g10797) );
  INVX0 U2030 ( .INP(g1861), .ZN(n1718) );
  NAND2X0 U2031 ( .IN1(g1845), .IN2(n1718), .QN(n1568) );
  NOR2X0 U2032 ( .IN1(g1864), .IN2(n1568), .QN(n1569) );
  INVX0 U2033 ( .INP(n1569), .ZN(n1375) );
  NAND2X0 U2034 ( .IN1(g1868), .IN2(n1375), .QN(n1376) );
  INVX0 U2035 ( .INP(n1903), .ZN(n1804) );
  NOR2X0 U2036 ( .IN1(n1733), .IN2(n1804), .QN(n1909) );
  NAND2X0 U2037 ( .IN1(n1376), .IN2(n1909), .QN(g6909) );
  INVX0 U2038 ( .INP(n1694), .ZN(n1961) );
  NAND2X0 U2039 ( .IN1(g627), .IN2(g643), .QN(n1664) );
  INVX0 U2040 ( .INP(n1664), .ZN(n1378) );
  INVX0 U2041 ( .INP(g646), .ZN(n1377) );
  NAND2X0 U2042 ( .IN1(n1378), .IN2(n1377), .QN(n1662) );
  NOR2X0 U2043 ( .IN1(g650), .IN2(n1662), .QN(n1590) );
  INVX0 U2044 ( .INP(n1590), .ZN(n1416) );
  INVX0 U2045 ( .INP(g654), .ZN(n1379) );
  INVX0 U2046 ( .INP(n1828), .ZN(n1603) );
  NOR2X0 U2047 ( .IN1(n1961), .IN2(n1603), .QN(n1663) );
  OR2X1 U2048 ( .IN1(g643), .IN2(g627), .Q(n1380) );
  NAND3X0 U2049 ( .IN1(n1663), .IN2(n1380), .IN3(n1664), .QN(g7441) );
  NAND2X0 U2050 ( .IN1(n1778), .IN2(n1942), .QN(n1826) );
  INVX0 U2051 ( .INP(n1826), .ZN(n1670) );
  OA21X1 U2052 ( .IN1(g611), .IN2(n1670), .IN3(n1940), .Q(n1005) );
  INVX0 U2053 ( .INP(n1005), .ZN(n1669) );
  AND2X1 U2054 ( .IN1(n1669), .IN2(g632), .Q(g4892) );
  AND2X1 U2055 ( .IN1(g1850), .IN2(n1727), .Q(g4904) );
  NAND2X0 U2056 ( .IN1(g18), .IN2(g213), .QN(n1629) );
  MUX21X1 U2057 ( .IN1(g1624), .IN2(n1629), .S(n2007), .Q(n1381) );
  INVX0 U2058 ( .INP(n1381), .ZN(g8773) );
  MUX21X1 U2059 ( .IN1(g1627), .IN2(n1696), .S(n2007), .Q(n1382) );
  INVX0 U2060 ( .INP(n1382), .ZN(g8774) );
  MUX21X1 U2061 ( .IN1(g1615), .IN2(n1495), .S(n2007), .Q(n1383) );
  INVX0 U2062 ( .INP(n1383), .ZN(g8770) );
  INVX0 U2063 ( .INP(g617), .ZN(n1941) );
  NOR2X0 U2064 ( .IN1(n1828), .IN2(n1941), .QN(n1771) );
  NAND2X0 U2065 ( .IN1(n1771), .IN2(n1945), .QN(n1384) );
  INVX0 U2066 ( .INP(n1384), .ZN(n2004) );
  AND2X1 U2067 ( .IN1(g736), .IN2(n2004), .Q(n1672) );
  NOR2X0 U2068 ( .IN1(n1961), .IN2(n1672), .QN(n1386) );
  NAND2X0 U2069 ( .IN1(g664), .IN2(n1384), .QN(n1385) );
  NAND2X0 U2070 ( .IN1(n1386), .IN2(n1385), .QN(g8649) );
  INVX0 U2071 ( .INP(g391), .ZN(n1387) );
  MUX21X1 U2072 ( .IN1(g391), .IN2(n1387), .S(g321), .Q(n1412) );
  INVX0 U2073 ( .INP(g401), .ZN(n1388) );
  MUX21X1 U2074 ( .IN1(g401), .IN2(n1388), .S(g327), .Q(n1411) );
  INVX0 U2075 ( .INP(g416), .ZN(n1396) );
  MUX21X1 U2076 ( .IN1(n1396), .IN2(g416), .S(g309), .Q(n1394) );
  INVX0 U2077 ( .INP(g421), .ZN(n1395) );
  MUX21X1 U2078 ( .IN1(n1395), .IN2(g421), .S(g312), .Q(n1393) );
  INVX0 U2079 ( .INP(g386), .ZN(n1389) );
  MUX21X1 U2080 ( .IN1(n1389), .IN2(g386), .S(g318), .Q(n1392) );
  INVX0 U2081 ( .INP(g396), .ZN(n1390) );
  MUX21X1 U2082 ( .IN1(n1390), .IN2(g396), .S(g324), .Q(n1391) );
  NAND4X0 U2083 ( .IN1(n1394), .IN2(n1393), .IN3(n1392), .IN4(n1391), .QN(
        n1410) );
  INVX0 U2084 ( .INP(g305), .ZN(n1460) );
  NOR2X0 U2085 ( .IN1(g435), .IN2(g431), .QN(n1401) );
  INVX0 U2086 ( .INP(g411), .ZN(n1403) );
  INVX0 U2087 ( .INP(g406), .ZN(n1402) );
  NAND4X0 U2088 ( .IN1(n1403), .IN2(n1402), .IN3(n1396), .IN4(n1395), .QN(
        n1399) );
  OR4X1 U2089 ( .IN1(g396), .IN2(g391), .IN3(g401), .IN4(g448), .Q(n1397) );
  OR4X1 U2090 ( .IN1(g426), .IN2(g386), .IN3(g452), .IN4(n1397), .Q(n1398) );
  OR4X1 U2091 ( .IN1(g444), .IN2(g440), .IN3(n1399), .IN4(n1398), .Q(n1400) );
  NAND4X0 U2092 ( .IN1(g374), .IN2(g382), .IN3(g369), .IN4(g378), .QN(n1459)
         );
  AO221X1 U2093 ( .IN1(g431), .IN2(g435), .IN3(n1401), .IN4(n1400), .IN5(n1459), .Q(n1461) );
  MUX21X1 U2094 ( .IN1(n1460), .IN2(g305), .S(n1461), .Q(n1408) );
  MUX21X1 U2095 ( .IN1(n1402), .IN2(g406), .S(g330), .Q(n1407) );
  MUX21X1 U2096 ( .IN1(n1403), .IN2(g411), .S(g333), .Q(n1406) );
  INVX0 U2097 ( .INP(g426), .ZN(n1404) );
  MUX21X1 U2098 ( .IN1(n1404), .IN2(g426), .S(g315), .Q(n1405) );
  NAND4X0 U2099 ( .IN1(n1408), .IN2(n1407), .IN3(n1406), .IN4(n1405), .QN(
        n1409) );
  NOR4X0 U2100 ( .IN1(n1412), .IN2(n1411), .IN3(n1410), .IN4(n1409), .QN(n1413) );
  NOR2X0 U2101 ( .IN1(n1413), .IN2(n1459), .QN(n1414) );
  NAND2X0 U2102 ( .IN1(n1414), .IN2(n1453), .QN(n1747) );
  INVX0 U2103 ( .INP(n1747), .ZN(g10788) );
  NAND2X0 U2104 ( .IN1(g654), .IN2(n1416), .QN(n1417) );
  NAND2X0 U2105 ( .IN1(n1417), .IN2(n1663), .QN(g7660) );
  INVX0 U2106 ( .INP(g1700), .ZN(n1008) );
  NAND2X0 U2107 ( .IN1(g109), .IN2(g757), .QN(n1744) );
  NAND2X0 U2108 ( .IN1(g878), .IN2(g876), .QN(n1743) );
  INVX0 U2109 ( .INP(n1419), .ZN(n1816) );
  NAND2X0 U2110 ( .IN1(n1816), .IN2(g881), .QN(n1422) );
  INVX0 U2111 ( .INP(n1420), .ZN(n1829) );
  NAND2X0 U2112 ( .IN1(n1829), .IN2(g877), .QN(n1421) );
  NAND2X0 U2113 ( .IN1(n1422), .IN2(n1421), .QN(n1423) );
  NOR2X0 U2114 ( .IN1(n1424), .IN2(n1423), .QN(g10515) );
  AND2X1 U2115 ( .IN1(g762), .IN2(g758), .Q(n1722) );
  NOR2X0 U2116 ( .IN1(g766), .IN2(n1722), .QN(n1426) );
  NAND3X0 U2117 ( .IN1(g762), .IN2(g758), .IN3(g766), .QN(n1544) );
  NOR2X0 U2118 ( .IN1(g590), .IN2(n1022), .QN(n1721) );
  NAND2X0 U2119 ( .IN1(n1544), .IN2(n1721), .QN(n1425) );
  NOR2X0 U2120 ( .IN1(n1426), .IN2(n1425), .QN(g5536) );
  INVX0 U2121 ( .INP(g770), .ZN(n1543) );
  NOR2X0 U2122 ( .IN1(n1544), .IN2(n1543), .QN(n1427) );
  NOR2X0 U2123 ( .IN1(g774), .IN2(n1427), .QN(n1429) );
  NAND2X0 U2124 ( .IN1(n1427), .IN2(g774), .QN(n1622) );
  NAND2X0 U2125 ( .IN1(n1622), .IN2(n1721), .QN(n1428) );
  NOR2X0 U2126 ( .IN1(n1429), .IN2(n1428), .QN(g6728) );
  NAND2X0 U2127 ( .IN1(g802), .IN2(g806), .QN(n1958) );
  NOR2X0 U2128 ( .IN1(n1957), .IN2(n1958), .QN(n1648) );
  NOR2X0 U2129 ( .IN1(n1648), .IN2(g810), .QN(n1431) );
  NAND2X0 U2130 ( .IN1(g810), .IN2(n1648), .QN(n1676) );
  NAND2X0 U2131 ( .IN1(n1676), .IN2(n1675), .QN(n1430) );
  NOR2X0 U2132 ( .IN1(n1431), .IN2(n1430), .QN(g6733) );
  INVX0 U2133 ( .INP(g1696), .ZN(n1699) );
  INVX0 U2134 ( .INP(n1881), .ZN(n1768) );
  NAND3X0 U2135 ( .IN1(g1766), .IN2(g1771), .IN3(g1776), .QN(n2014) );
  NOR2X0 U2136 ( .IN1(n1768), .IN2(n2014), .QN(n1482) );
  NOR2X0 U2137 ( .IN1(n1482), .IN2(g1781), .QN(n1433) );
  NAND2X0 U2138 ( .IN1(g1781), .IN2(n1482), .QN(n1571) );
  NAND2X0 U2139 ( .IN1(n1571), .IN2(n1636), .QN(n1432) );
  NOR2X0 U2140 ( .IN1(n1433), .IN2(n1432), .QN(g6516) );
  NAND2X0 U2141 ( .IN1(g1786), .IN2(g1791), .QN(n1434) );
  NOR2X0 U2142 ( .IN1(n2014), .IN2(n1434), .QN(n1435) );
  NAND2X0 U2143 ( .IN1(g1781), .IN2(n1435), .QN(n1572) );
  NOR2X0 U2144 ( .IN1(n1768), .IN2(n1572), .QN(n1570) );
  NOR2X0 U2145 ( .IN1(n1570), .IN2(g1796), .QN(n1437) );
  NAND2X0 U2146 ( .IN1(g1796), .IN2(n1570), .QN(n1479) );
  NAND2X0 U2147 ( .IN1(n1479), .IN2(n1636), .QN(n1436) );
  NOR2X0 U2148 ( .IN1(n1437), .IN2(n1436), .QN(g7541) );
  INVX0 U2149 ( .INP(g778), .ZN(n1621) );
  NOR2X0 U2150 ( .IN1(n1622), .IN2(n1621), .QN(n1438) );
  NOR2X0 U2151 ( .IN1(g782), .IN2(n1438), .QN(n1440) );
  NAND2X0 U2152 ( .IN1(n1438), .IN2(g782), .QN(n1627) );
  NAND2X0 U2153 ( .IN1(n1627), .IN2(n1721), .QN(n1439) );
  NOR2X0 U2154 ( .IN1(n1440), .IN2(n1439), .QN(g7705) );
  INVX0 U2155 ( .INP(g814), .ZN(n1677) );
  NOR2X0 U2156 ( .IN1(n1677), .IN2(n1676), .QN(n1441) );
  NOR2X0 U2157 ( .IN1(n1441), .IN2(g818), .QN(n1443) );
  NAND2X0 U2158 ( .IN1(g818), .IN2(n1441), .QN(n1594) );
  NAND2X0 U2159 ( .IN1(n1594), .IN2(n1675), .QN(n1442) );
  NOR2X0 U2160 ( .IN1(n1443), .IN2(n1442), .QN(g7709) );
  NOR2X0 U2161 ( .IN1(g1218), .IN2(n1289), .QN(n1445) );
  NAND3X0 U2162 ( .IN1(g1218), .IN2(n1289), .IN3(n1763), .QN(n1514) );
  NOR2X0 U2163 ( .IN1(g1212), .IN2(n1022), .QN(n1560) );
  NAND2X0 U2164 ( .IN1(n1514), .IN2(n1560), .QN(n1444) );
  NOR2X0 U2165 ( .IN1(n1445), .IN2(n1444), .QN(g7632) );
  INVX0 U2166 ( .INP(g786), .ZN(n1626) );
  NOR2X0 U2167 ( .IN1(n1627), .IN2(n1626), .QN(n1446) );
  NOR2X0 U2168 ( .IN1(g790), .IN2(n1446), .QN(n1448) );
  NAND2X0 U2169 ( .IN1(n1446), .IN2(g790), .QN(n2011) );
  NAND2X0 U2170 ( .IN1(n2011), .IN2(n1721), .QN(n1447) );
  NOR2X0 U2171 ( .IN1(n1448), .IN2(n1447), .QN(g8244) );
  INVX0 U2172 ( .INP(g1223), .ZN(n1515) );
  NOR2X0 U2173 ( .IN1(n1515), .IN2(n1514), .QN(n1449) );
  NOR2X0 U2174 ( .IN1(n1449), .IN2(g1227), .QN(n1452) );
  INVX0 U2175 ( .INP(n1514), .ZN(n1450) );
  NAND3X0 U2176 ( .IN1(g1227), .IN2(g1223), .IN3(n1450), .QN(n1559) );
  NAND2X0 U2177 ( .IN1(n1559), .IN2(n1560), .QN(n1451) );
  NOR2X0 U2178 ( .IN1(n1452), .IN2(n1451), .QN(g7586) );
  NOR2X0 U2179 ( .IN1(n1467), .IN2(g369), .QN(n1455) );
  NOR2X0 U2180 ( .IN1(g869), .IN2(n1022), .QN(n1527) );
  NAND2X0 U2181 ( .IN1(n1483), .IN2(n1527), .QN(n1454) );
  NOR2X0 U2182 ( .IN1(n1455), .IN2(n1454), .QN(g11320) );
  NBUFFX2 U2183 ( .INP(n1470), .Z(n1964) );
  MUX21X1 U2184 ( .IN1(g501), .IN2(g506), .S(n1964), .Q(g11335) );
  NBUFFX2 U2185 ( .INP(n1470), .Z(n1968) );
  MUX21X1 U2186 ( .IN1(g516), .IN2(g476), .S(n1968), .Q(g11338) );
  MUX21X1 U2187 ( .IN1(g421), .IN2(g452), .S(n1968), .Q(g11257) );
  MUX21X1 U2188 ( .IN1(g406), .IN2(g411), .S(n1968), .Q(g11268) );
  INVX0 U2189 ( .INP(g374), .ZN(n1484) );
  NOR2X0 U2190 ( .IN1(n1484), .IN2(n1483), .QN(n1456) );
  NOR2X0 U2191 ( .IN1(n1456), .IN2(g378), .QN(n1458) );
  NAND2X0 U2192 ( .IN1(g378), .IN2(n1456), .QN(n1526) );
  NAND2X0 U2193 ( .IN1(n1526), .IN2(n1527), .QN(n1457) );
  NOR2X0 U2194 ( .IN1(n1458), .IN2(n1457), .QN(g11291) );
  MUX21X1 U2195 ( .IN1(g411), .IN2(g416), .S(n1968), .Q(g11269) );
  NAND2X0 U2196 ( .IN1(n1460), .IN2(n1459), .QN(n1462) );
  NAND2X0 U2197 ( .IN1(n1462), .IN2(n1461), .QN(n1463) );
  MUX21X1 U2198 ( .IN1(n1463), .IN2(g426), .S(n1964), .Q(g11256) );
  NOR2X0 U2199 ( .IN1(g10788), .IN2(g971), .QN(n1466) );
  NAND2X0 U2200 ( .IN1(g971), .IN2(g10788), .QN(n1610) );
  NAND2X0 U2201 ( .IN1(g869), .IN2(n1743), .QN(n1464) );
  OA21X1 U2202 ( .IN1(g757), .IN2(n1464), .IN3(g109), .Q(n1609) );
  NAND2X0 U2203 ( .IN1(n1610), .IN2(n1609), .QN(n1465) );
  NOR2X0 U2204 ( .IN1(n1466), .IN2(n1465), .QN(g11349) );
  NOR2X0 U2205 ( .IN1(n1467), .IN2(g456), .QN(n1473) );
  NOR2X0 U2206 ( .IN1(n1562), .IN2(n1468), .QN(n1471) );
  NOR2X0 U2207 ( .IN1(g868), .IN2(n1022), .QN(n1728) );
  NAND2X0 U2208 ( .IN1(n1511), .IN2(n1728), .QN(n1472) );
  NOR2X0 U2209 ( .IN1(n1473), .IN2(n1472), .QN(g11340) );
  NOR2X0 U2210 ( .IN1(g11561), .IN2(g1336), .QN(n1476) );
  NAND3X0 U2211 ( .IN1(g109), .IN2(g1206), .IN3(g1361), .QN(n2023) );
  NAND2X0 U2212 ( .IN1(g1212), .IN2(n2023), .QN(n1474) );
  OA21X1 U2213 ( .IN1(g108), .IN2(n1474), .IN3(g109), .Q(n1519) );
  NAND2X0 U2214 ( .IN1(n1521), .IN2(n1519), .QN(n1475) );
  NOR2X0 U2215 ( .IN1(n1476), .IN2(n1475), .QN(g11636) );
  AND2X1 U2216 ( .IN1(g1690), .IN2(g1687), .Q(g6955) );
  NAND3X0 U2218 ( .IN1(g1336), .IN2(n1519), .IN3(g11561), .QN(n1477) );
  NOR2X0 U2219 ( .IN1(n1507), .IN2(n1477), .QN(n1524) );
  OA21X1 U2220 ( .IN1(n1507), .IN2(n1521), .IN3(n1519), .Q(n1478) );
  NBUFFX2 U2221 ( .INP(g1346), .Z(n1525) );
  MUX21X1 U2222 ( .IN1(n1524), .IN2(n1478), .S(n1525), .Q(g11640) );
  INVX0 U2225 ( .INP(g1801), .ZN(n2019) );
  NOR2X0 U2226 ( .IN1(n2019), .IN2(n1479), .QN(n1639) );
  INVX0 U2227 ( .INP(n1639), .ZN(n1637) );
  NAND2X0 U2228 ( .IN1(n2019), .IN2(n1479), .QN(n1480) );
  AND3X1 U2229 ( .IN1(n1636), .IN2(n1637), .IN3(n1480), .Q(g7930) );
  AND3X1 U2230 ( .IN1(g1766), .IN2(g1771), .IN3(n1881), .Q(n1619) );
  NOR2X0 U2231 ( .IN1(g1776), .IN2(n1619), .QN(n1481) );
  NOR3X0 U2232 ( .IN1(g1713), .IN2(n1482), .IN3(n1481), .QN(g6508) );
  INVX0 U2233 ( .INP(n1483), .ZN(n1485) );
  OA221X1 U2234 ( .IN1(g374), .IN2(n1485), .IN3(n1484), .IN4(n1483), .IN5(
        n1527), .Q(g11290) );
  AND2X1 U2235 ( .IN1(g109), .IN2(g213), .Q(g6829) );
  INVX0 U2236 ( .INP(g18), .ZN(n1606) );
  NOR3X0 U2237 ( .IN1(g1840), .IN2(n1591), .IN3(n1487), .QN(n1540) );
  INVX0 U2238 ( .INP(n1540), .ZN(n1739) );
  NAND2X0 U2239 ( .IN1(g1822), .IN2(n1487), .QN(n1791) );
  NAND3X0 U2240 ( .IN1(n1739), .IN2(n1791), .IN3(n1592), .QN(n1492) );
  INVX0 U2241 ( .INP(g1891), .ZN(n2000) );
  NAND3X0 U2242 ( .IN1(n1487), .IN2(n1486), .IN3(g1828), .QN(n1798) );
  OA21X1 U2243 ( .IN1(g1828), .IN2(n1791), .IN3(n1798), .Q(n1503) );
  NAND2X0 U2244 ( .IN1(n1503), .IN2(n1592), .QN(n1784) );
  NAND3X0 U2245 ( .IN1(g1882), .IN2(g1872), .IN3(n1784), .QN(n1995) );
  NOR2X0 U2246 ( .IN1(n2000), .IN2(n1995), .QN(n1753) );
  NAND3X0 U2247 ( .IN1(g1900), .IN2(g1909), .IN3(g1918), .QN(n1756) );
  INVX0 U2248 ( .INP(n1756), .ZN(n1488) );
  AND3X1 U2249 ( .IN1(n1753), .IN2(g1927), .IN3(n1488), .Q(n1973) );
  NAND2X0 U2250 ( .IN1(g1936), .IN2(n1973), .QN(n1735) );
  INVX0 U2251 ( .INP(g1945), .ZN(n1738) );
  INVX0 U2252 ( .INP(g1882), .ZN(n1490) );
  INVX0 U2253 ( .INP(g1872), .ZN(n1489) );
  NAND2X0 U2254 ( .IN1(n1490), .IN2(n1489), .QN(n1491) );
  NOR2X0 U2255 ( .IN1(n1784), .IN2(n1491), .QN(n1993) );
  NAND2X0 U2256 ( .IN1(n1993), .IN2(n2000), .QN(n1754) );
  INVX0 U2257 ( .INP(g1900), .ZN(n1848) );
  INVX0 U2258 ( .INP(g1909), .ZN(n1824) );
  INVX0 U2259 ( .INP(g1918), .ZN(n1932) );
  NAND3X0 U2260 ( .IN1(n1848), .IN2(n1824), .IN3(n1932), .QN(n1755) );
  NOR3X0 U2261 ( .IN1(g1927), .IN2(n1754), .IN3(n1755), .QN(n1972) );
  INVX0 U2262 ( .INP(g1936), .ZN(n1976) );
  NAND2X0 U2263 ( .IN1(n1972), .IN2(n1976), .QN(n1734) );
  INVX0 U2264 ( .INP(g1857), .ZN(n1908) );
  INVX0 U2265 ( .INP(n1733), .ZN(n1891) );
  AO221X1 U2266 ( .IN1(n1739), .IN2(n1892), .IN3(n1739), .IN4(n1908), .IN5(
        n1891), .Q(n1749) );
  AO221X1 U2267 ( .IN1(g1945), .IN2(n1735), .IN3(n1738), .IN4(n1734), .IN5(
        n1749), .Q(n1564) );
  INVX0 U2268 ( .INP(n1564), .ZN(n1732) );
  NAND2X0 U2269 ( .IN1(n1492), .IN2(n1732), .QN(n1493) );
  NOR2X0 U2270 ( .IN1(n1606), .IN2(n1494), .QN(g9266) );
  AND2X1 U2271 ( .IN1(g109), .IN2(g243), .Q(g6819) );
  INVX0 U2272 ( .INP(g1428), .ZN(n1496) );
  MUX21X1 U2273 ( .IN1(g1428), .IN2(n1496), .S(n1495), .Q(n1497) );
  NOR2X0 U2274 ( .IN1(n1022), .IN2(n1497), .QN(g8769) );
  AND2X1 U2275 ( .IN1(g109), .IN2(g1377), .Q(g6828) );
  AND2X1 U2276 ( .IN1(g109), .IN2(g1380), .Q(g6830) );
  INVX0 U2277 ( .INP(g1432), .ZN(n1577) );
  MUX21X1 U2278 ( .IN1(g1432), .IN2(n1577), .S(n1629), .Q(n1498) );
  NOR2X0 U2279 ( .IN1(n1022), .IN2(n1498), .QN(g8765) );
  AND2X1 U2280 ( .IN1(g109), .IN2(g1499), .Q(g6198) );
  NOR2X0 U2281 ( .IN1(g1393), .IN2(g1394), .QN(n1499) );
  NOR3X0 U2282 ( .IN1(n1499), .IN2(g115), .IN3(n1022), .QN(g6747) );
  AND2X1 U2283 ( .IN1(g1849), .IN2(n1727), .Q(g4903) );
  INVX0 U2284 ( .INP(g822), .ZN(n1595) );
  NOR2X0 U2285 ( .IN1(n1595), .IN2(n1594), .QN(n1501) );
  INVX0 U2286 ( .INP(g826), .ZN(n1500) );
  INVX0 U2287 ( .INP(n1501), .ZN(n1597) );
  OA221X1 U2288 ( .IN1(g826), .IN2(n1501), .IN3(n1500), .IN4(n1597), .IN5(
        n1675), .Q(g8245) );
  NOR2X0 U2289 ( .IN1(n1487), .IN2(n1788), .QN(n1790) );
  NAND2X0 U2290 ( .IN1(n1790), .IN2(g1822), .QN(n1502) );
  AO21X1 U2291 ( .IN1(n1503), .IN2(n1502), .IN3(n1564), .Q(n1504) );
  NAND2X0 U2292 ( .IN1(n1788), .IN2(n1504), .QN(n1505) );
  OA221X1 U2293 ( .IN1(n1505), .IN2(n1804), .IN3(n1788), .IN4(n1504), .IN5(g18), .Q(g9272) );
  AND2X1 U2294 ( .IN1(g109), .IN2(g237), .Q(g6821) );
  INVX0 U2295 ( .INP(g1444), .ZN(n1580) );
  NAND2X0 U2296 ( .IN1(g18), .IN2(g231), .QN(n1565) );
  INVX0 U2297 ( .INP(n1565), .ZN(n1862) );
  MUX21X1 U2298 ( .IN1(n1580), .IN2(g1444), .S(n1862), .Q(n1506) );
  NOR2X0 U2299 ( .IN1(n1022), .IN2(n1506), .QN(g8768) );
  INVX0 U2300 ( .INP(n1521), .ZN(n1508) );
  OA221X1 U2301 ( .IN1(g1341), .IN2(n1508), .IN3(n1507), .IN4(n1521), .IN5(
        n1519), .Q(g11639) );
  AND2X1 U2302 ( .IN1(g109), .IN2(g1400), .Q(g6841) );
  INVX0 U2303 ( .INP(n1610), .ZN(n1509) );
  INVX0 U2304 ( .INP(g976), .ZN(n1611) );
  OA221X1 U2305 ( .IN1(g976), .IN2(n1509), .IN3(n1611), .IN4(n1610), .IN5(
        n1609), .Q(g11391) );
  INVX0 U2306 ( .INP(n1957), .ZN(n1510) );
  INVX0 U2307 ( .INP(g802), .ZN(n1646) );
  OA221X1 U2308 ( .IN1(n1510), .IN2(g802), .IN3(n1957), .IN4(n1646), .IN5(
        n1675), .Q(g5543) );
  NOR2X0 U2309 ( .IN1(n1512), .IN2(n1511), .QN(n1731) );
  INVX0 U2310 ( .INP(n1731), .ZN(n1729) );
  NAND2X0 U2311 ( .IN1(n1512), .IN2(n1511), .QN(n1513) );
  AND3X1 U2312 ( .IN1(n1729), .IN2(n1728), .IN3(n1513), .Q(g11372) );
  AND2X1 U2313 ( .IN1(g109), .IN2(g1368), .Q(g6823) );
  INVX0 U2314 ( .INP(g1419), .ZN(n1578) );
  NOR2X0 U2315 ( .IN1(n1022), .IN2(n1578), .QN(g6193) );
  AND2X1 U2316 ( .IN1(n1289), .IN2(g1218), .Q(n1516) );
  OA221X1 U2317 ( .IN1(g1223), .IN2(n1516), .IN3(n1515), .IN4(n1514), .IN5(
        n1560), .Q(g7581) );
  AND2X1 U2318 ( .IN1(g109), .IN2(g1365), .Q(g6834) );
  AND2X1 U2319 ( .IN1(g109), .IN2(g1453), .Q(g6180) );
  NOR2X0 U2320 ( .IN1(g1453), .IN2(n1022), .QN(n1518) );
  INVX0 U2321 ( .INP(g1494), .ZN(n1660) );
  XNOR3X1 U2322 ( .IN1(g1508), .IN2(g1499), .IN3(n1660), .Q(n1517) );
  MUX21X1 U2323 ( .IN1(g6180), .IN2(n1518), .S(n1517), .Q(g5770) );
  INVX0 U2324 ( .INP(g1351), .ZN(n1523) );
  NAND2X0 U2325 ( .IN1(g1341), .IN2(n1525), .QN(n1520) );
  OA21X1 U2326 ( .IN1(n1521), .IN2(n1520), .IN3(n1519), .Q(n1522) );
  OA222X1 U2327 ( .IN1(g1351), .IN2(n1525), .IN3(g1351), .IN4(n1524), .IN5(
        n1523), .IN6(n1522), .Q(g11641) );
  AND4X1 U2328 ( .IN1(g1351), .IN2(g1336), .IN3(g1341), .IN4(n1525), .Q(g4114)
         );
  INVX0 U2329 ( .INP(n1526), .ZN(n1528) );
  OA21X1 U2330 ( .IN1(g382), .IN2(n1528), .IN3(n1527), .Q(g11292) );
  AND2X1 U2331 ( .IN1(g109), .IN2(g178), .Q(g6786) );
  INVX0 U2332 ( .INP(g174), .ZN(n1617) );
  NOR4X0 U2333 ( .IN1(g119), .IN2(g158), .IN3(g131), .IN4(n1617), .QN(n1533)
         );
  INVX0 U2334 ( .INP(g127), .ZN(n1539) );
  INVX0 U2335 ( .INP(g139), .ZN(n1716) );
  NAND4X0 U2336 ( .IN1(g182), .IN2(g170), .IN3(n1539), .IN4(n1716), .QN(n1531)
         );
  OR4X1 U2337 ( .IN1(g148), .IN2(g143), .IN3(g162), .IN4(g153), .Q(n1530) );
  NAND4X0 U2338 ( .IN1(g18), .IN2(g115), .IN3(g166), .IN4(g6786), .QN(n1529)
         );
  NOR4X0 U2339 ( .IN1(g135), .IN2(n1531), .IN3(n1530), .IN4(n1529), .QN(n1532)
         );
  AO22X1 U2340 ( .IN1(g109), .IN2(g123), .IN3(n1533), .IN4(n1532), .Q(g7032)
         );
  INVX0 U2341 ( .INP(n1571), .ZN(n1534) );
  INVX0 U2342 ( .INP(g1786), .ZN(n2016) );
  OA221X1 U2343 ( .IN1(g1786), .IN2(n1534), .IN3(n2016), .IN4(n1571), .IN5(
        n1636), .Q(g6525) );
  INVX0 U2344 ( .INP(g1482), .ZN(n1536) );
  OA221X1 U2345 ( .IN1(n1537), .IN2(n1536), .IN3(n1535), .IN4(g1482), .IN5(
        g109), .Q(g8046) );
  MUX21X1 U2346 ( .IN1(g566), .IN2(g231), .S(g18), .Q(g6035) );
  INVX0 U2347 ( .INP(g6035), .ZN(n1538) );
  OA221X1 U2348 ( .IN1(g127), .IN2(g6035), .IN3(n1539), .IN4(n1538), .IN5(g109), .Q(g8047) );
  OA221X1 U2349 ( .IN1(g1840), .IN2(n1540), .IN3(g1840), .IN4(n1564), .IN5(
        n1733), .Q(n1541) );
  MUX21X1 U2350 ( .IN1(n1591), .IN2(g1834), .S(n1541), .Q(n1542) );
  NOR2X0 U2351 ( .IN1(n1606), .IN2(n1542), .QN(g9555) );
  AND2X1 U2352 ( .IN1(g109), .IN2(g1383), .Q(g6832) );
  INVX0 U2353 ( .INP(n1544), .ZN(n1545) );
  OA221X1 U2354 ( .IN1(n1545), .IN2(g770), .IN3(n1544), .IN4(n1543), .IN5(
        n1721), .Q(g6123) );
  AND2X1 U2355 ( .IN1(g109), .IN2(g1389), .Q(g6334) );
  NOR2X0 U2356 ( .IN1(n1022), .IN2(g1389), .QN(n1555) );
  NOR4X0 U2357 ( .IN1(g1389), .IN2(g1386), .IN3(g1397), .IN4(g1383), .QN(n1552) );
  NOR4X0 U2358 ( .IN1(g219), .IN2(g213), .IN3(g186), .IN4(g248), .QN(n1551) );
  NOR3X0 U2359 ( .IN1(g237), .IN2(g207), .IN3(g1380), .QN(n1550) );
  NOR4X0 U2360 ( .IN1(g1400), .IN2(g1365), .IN3(g1368), .IN4(g1377), .QN(n1548) );
  NOR4X0 U2361 ( .IN1(g197), .IN2(g1371), .IN3(g1362), .IN4(g1374), .QN(n1547)
         );
  NOR4X0 U2362 ( .IN1(g231), .IN2(g225), .IN3(g192), .IN4(g243), .QN(n1546) );
  AND3X1 U2363 ( .IN1(n1548), .IN2(n1547), .IN3(n1546), .Q(n1549) );
  NAND4X0 U2364 ( .IN1(n1552), .IN2(n1551), .IN3(n1550), .IN4(n1549), .QN(
        n1558) );
  NAND2X0 U2365 ( .IN1(n1558), .IN2(g201), .QN(n1553) );
  XNOR3X1 U2366 ( .IN1(g197), .IN2(g1386), .IN3(n1553), .Q(n1554) );
  MUX21X1 U2367 ( .IN1(n1555), .IN2(g6334), .S(n1554), .Q(g5755) );
  INVX0 U2368 ( .INP(n1556), .ZN(n1633) );
  OA21X1 U2369 ( .IN1(g12), .IN2(n1633), .IN3(g109), .Q(g5445) );
  AND2X1 U2370 ( .IN1(g109), .IN2(g1397), .Q(g6839) );
  AND2X1 U2371 ( .IN1(n1669), .IN2(g630), .Q(g4890) );
  NOR2X0 U2372 ( .IN1(n1022), .IN2(g201), .QN(g6331) );
  INVX0 U2373 ( .INP(g6331), .ZN(n1557) );
  NOR2X0 U2374 ( .IN1(n1558), .IN2(n1557), .QN(g6163) );
  AND2X1 U2375 ( .IN1(g6163), .IN2(g1394), .Q(g6179) );
  INVX0 U2376 ( .INP(n1559), .ZN(n1561) );
  OA21X1 U2377 ( .IN1(g1231), .IN2(n1561), .IN3(n1560), .Q(g7590) );
  AND3X1 U2378 ( .IN1(g109), .IN2(g741), .IN3(g742), .Q(g3407) );
  NOR2X0 U2379 ( .IN1(n1964), .IN2(n1562), .QN(n1563) );
  OA21X1 U2380 ( .IN1(g471), .IN2(n1563), .IN3(n1728), .Q(g11380) );
  AND2X1 U2381 ( .IN1(g109), .IN2(g1374), .Q(g6332) );
  OA221X1 U2382 ( .IN1(n1732), .IN2(g1822), .IN3(n1564), .IN4(g1828), .IN5(g18), .Q(g9269) );
  OA21X1 U2383 ( .IN1(g9), .IN2(n1633), .IN3(g109), .Q(g5421) );
  OA21X1 U2384 ( .IN1(g18), .IN2(g1627), .IN3(n1565), .Q(n1567) );
  INVX0 U2385 ( .INP(g1474), .ZN(n1566) );
  INVX0 U2386 ( .INP(n1567), .ZN(n1781) );
  OA221X1 U2387 ( .IN1(n1567), .IN2(n1566), .IN3(n1781), .IN4(g1474), .IN5(
        g109), .Q(g8040) );
  AND2X1 U2388 ( .IN1(g109), .IN2(g192), .Q(g6838) );
  OA221X1 U2389 ( .IN1(n1569), .IN2(g1864), .IN3(n1569), .IN4(n1568), .IN5(
        n1909), .Q(g6795) );
  AND3X1 U2390 ( .IN1(g109), .IN2(g743), .IN3(g744), .Q(g3418) );
  INVX0 U2391 ( .INP(g1515), .ZN(n1579) );
  NOR2X0 U2392 ( .IN1(n1022), .IN2(n1579), .QN(g6205) );
  INVX0 U2393 ( .INP(g1791), .ZN(n2015) );
  NOR2X0 U2394 ( .IN1(n1570), .IN2(n2015), .QN(n1574) );
  NOR2X0 U2395 ( .IN1(n2016), .IN2(n1571), .QN(n1573) );
  OA221X1 U2396 ( .IN1(n1574), .IN2(n1573), .IN3(n1574), .IN4(n1572), .IN5(
        n1636), .Q(g6983) );
  MUX21X1 U2397 ( .IN1(g563), .IN2(g225), .S(g18), .Q(g6026) );
  INVX0 U2398 ( .INP(g170), .ZN(n1576) );
  INVX0 U2399 ( .INP(g6026), .ZN(n1575) );
  OA221X1 U2400 ( .IN1(g170), .IN2(g6026), .IN3(n1576), .IN4(n1575), .IN5(g109), .Q(g8050) );
  AND2X1 U2401 ( .IN1(g109), .IN2(g1520), .Q(g6224) );
  INVX0 U2402 ( .INP(g1440), .ZN(n1667) );
  NOR4X0 U2403 ( .IN1(n1579), .IN2(n1578), .IN3(n1577), .IN4(n1667), .QN(n1585) );
  NAND2X0 U2404 ( .IN1(g1428), .IN2(g1424), .QN(n1583) );
  INVX0 U2405 ( .INP(g1448), .ZN(n1631) );
  NOR4X0 U2406 ( .IN1(g1403), .IN2(g1411), .IN3(n1580), .IN4(n1631), .QN(n1581) );
  NAND4X0 U2407 ( .IN1(g1436), .IN2(n1581), .IN3(n1710), .IN4(g6224), .QN(
        n1582) );
  NOR4X0 U2408 ( .IN1(g1415), .IN2(g1407), .IN3(n1583), .IN4(n1582), .QN(n1584) );
  AO22X1 U2409 ( .IN1(g109), .IN2(g1), .IN3(n1585), .IN4(n1584), .Q(g6679) );
  AND2X1 U2410 ( .IN1(g109), .IN2(g1424), .Q(g6234) );
  AND2X1 U2411 ( .IN1(g109), .IN2(g207), .Q(g6831) );
  NOR2X0 U2412 ( .IN1(n1611), .IN2(n1586), .QN(n1613) );
  INVX0 U2413 ( .INP(g986), .ZN(n1589) );
  NAND2X0 U2414 ( .IN1(g976), .IN2(g981), .QN(n1587) );
  OA21X1 U2415 ( .IN1(n1610), .IN2(n1587), .IN3(n1609), .Q(n1588) );
  OA222X1 U2416 ( .IN1(g986), .IN2(g981), .IN3(g986), .IN4(n1613), .IN5(n1589), 
        .IN6(n1588), .Q(g11393) );
  AND4X1 U2417 ( .IN1(g986), .IN2(g971), .IN3(g976), .IN4(g981), .Q(g3506) );
  OA221X1 U2418 ( .IN1(n1590), .IN2(g650), .IN3(n1590), .IN4(n1662), .IN5(
        n1663), .Q(g7137) );
  INVX0 U2419 ( .INP(n1851), .ZN(n1915) );
  NAND2X0 U2420 ( .IN1(g1950), .IN2(n1915), .QN(n1853) );
  NOR4X0 U2421 ( .IN1(g1834), .IN2(g1828), .IN3(g1840), .IN4(n1592), .QN(n1795) );
  AO21X1 U2422 ( .IN1(n1733), .IN2(n1795), .IN3(g1840), .Q(n1593) );
  AND3X1 U2423 ( .IN1(g18), .IN2(n1853), .IN3(n1593), .Q(g8384) );
  AND2X1 U2424 ( .IN1(g109), .IN2(g148), .Q(g6759) );
  NAND2X0 U2425 ( .IN1(n1595), .IN2(n1594), .QN(n1596) );
  AND3X1 U2426 ( .IN1(n1597), .IN2(n1675), .IN3(n1596), .Q(g8024) );
  AND2X1 U2427 ( .IN1(g109), .IN2(g186), .Q(g6833) );
  OA21X1 U2428 ( .IN1(g591), .IN2(g605), .IN3(g599), .Q(n1805) );
  NOR2X0 U2429 ( .IN1(g677), .IN2(g668), .QN(n1599) );
  NOR4X0 U2430 ( .IN1(g686), .IN2(g695), .IN3(g658), .IN4(g713), .QN(n1598) );
  INVX0 U2431 ( .INP(g704), .ZN(n1921) );
  NAND4X0 U2432 ( .IN1(n1805), .IN2(n1599), .IN3(n1598), .IN4(n1921), .QN(
        n1772) );
  NOR2X0 U2433 ( .IN1(g722), .IN2(n1772), .QN(n1868) );
  INVX0 U2434 ( .INP(g731), .ZN(n1873) );
  INVX0 U2435 ( .INP(g722), .ZN(n1777) );
  NAND2X0 U2436 ( .IN1(g677), .IN2(g668), .QN(n1811) );
  NAND3X0 U2437 ( .IN1(g704), .IN2(g686), .IN3(g695), .QN(n1917) );
  NOR2X0 U2438 ( .IN1(n1811), .IN2(n1917), .QN(n1600) );
  INVX0 U2439 ( .INP(n1805), .ZN(n1810) );
  NAND4X0 U2440 ( .IN1(g658), .IN2(g713), .IN3(n1600), .IN4(n1810), .QN(n1773)
         );
  NOR2X0 U2441 ( .IN1(n1777), .IN2(n1773), .QN(n1869) );
  NAND3X0 U2442 ( .IN1(g611), .IN2(g591), .IN3(n1941), .QN(n1693) );
  INVX0 U2443 ( .INP(n1693), .ZN(n1601) );
  OA221X1 U2444 ( .IN1(n1601), .IN2(g639), .IN3(n1601), .IN4(n1826), .IN5(
        n1603), .Q(n1774) );
  OA221X1 U2445 ( .IN1(g731), .IN2(n1868), .IN3(n1873), .IN4(n1869), .IN5(
        n1774), .Q(n1726) );
  NOR2X0 U2446 ( .IN1(n1726), .IN2(n1693), .QN(n1602) );
  NAND2X0 U2447 ( .IN1(n1601), .IN2(n1726), .QN(n1687) );
  NOR2X0 U2448 ( .IN1(g622), .IN2(n1687), .QN(n1705) );
  AO221X1 U2449 ( .IN1(n1603), .IN2(g617), .IN3(n1603), .IN4(n1602), .IN5(
        n1705), .Q(n1604) );
  MUX21X1 U2450 ( .IN1(n1945), .IN2(g611), .S(n1604), .Q(n1605) );
  NOR2X0 U2451 ( .IN1(n1606), .IN2(n1605), .QN(g9721) );
  MUX21X1 U2452 ( .IN1(g569), .IN2(g237), .S(g18), .Q(g6038) );
  INVX0 U2453 ( .INP(g131), .ZN(n1608) );
  INVX0 U2454 ( .INP(g6038), .ZN(n1607) );
  OA221X1 U2455 ( .IN1(g131), .IN2(g6038), .IN3(n1608), .IN4(n1607), .IN5(g109), .Q(g8044) );
  OA21X1 U2456 ( .IN1(n1611), .IN2(n1610), .IN3(n1609), .Q(n1612) );
  NAND2X0 U2457 ( .IN1(g18), .IN2(g192), .QN(n1615) );
  INVX0 U2458 ( .INP(g1458), .ZN(n1614) );
  INVX0 U2459 ( .INP(n1615), .ZN(n1840) );
  OA221X1 U2460 ( .IN1(n1615), .IN2(n1614), .IN3(n1840), .IN4(g1458), .IN5(
        g109), .Q(g8042) );
  MUX21X1 U2461 ( .IN1(g560), .IN2(g219), .S(g18), .Q(g6015) );
  INVX0 U2462 ( .INP(g6015), .ZN(n1616) );
  OA221X1 U2463 ( .IN1(g174), .IN2(g6015), .IN3(n1617), .IN4(n1616), .IN5(g109), .Q(g8054) );
  INVX0 U2464 ( .INP(g1766), .ZN(n1767) );
  NOR2X0 U2465 ( .IN1(n1767), .IN2(n1768), .QN(n1618) );
  NOR2X0 U2466 ( .IN1(g1771), .IN2(n1618), .QN(n1620) );
  NOR3X0 U2467 ( .IN1(n1620), .IN2(g1713), .IN3(n1619), .QN(g6502) );
  AND2X1 U2468 ( .IN1(g109), .IN2(g1407), .Q(g6216) );
  AND2X1 U2469 ( .IN1(g109), .IN2(g225), .Q(g6826) );
  INVX0 U2470 ( .INP(n1622), .ZN(n1623) );
  OA221X1 U2471 ( .IN1(n1623), .IN2(g778), .IN3(n1622), .IN4(n1621), .IN5(
        n1721), .Q(g7191) );
  AND2X1 U2472 ( .IN1(g109), .IN2(g219), .Q(g6827) );
  AND2X1 U2473 ( .IN1(g109), .IN2(g197), .Q(g6333) );
  MUX21X1 U2474 ( .IN1(g549), .IN2(g192), .S(g18), .Q(g6049) );
  INVX0 U2475 ( .INP(g166), .ZN(n1625) );
  INVX0 U2476 ( .INP(g6049), .ZN(n1624) );
  OA221X1 U2477 ( .IN1(g166), .IN2(g6049), .IN3(n1625), .IN4(n1624), .IN5(g109), .Q(g8049) );
  INVX0 U2478 ( .INP(n1627), .ZN(n1628) );
  OA221X1 U2479 ( .IN1(n1628), .IN2(g786), .IN3(n1627), .IN4(n1626), .IN5(
        n1721), .Q(g8019) );
  OA21X1 U2480 ( .IN1(g18), .IN2(g1615), .IN3(n1629), .Q(n1630) );
  INVX0 U2481 ( .INP(g1486), .ZN(n1708) );
  INVX0 U2482 ( .INP(n1630), .ZN(n1818) );
  OA221X1 U2483 ( .IN1(n1630), .IN2(n1708), .IN3(n1818), .IN4(g1486), .IN5(
        g109), .Q(g8052) );
  AND2X1 U2484 ( .IN1(g18), .IN2(g237), .Q(n1969) );
  MUX21X1 U2485 ( .IN1(n1631), .IN2(g1448), .S(n1969), .Q(n1632) );
  NOR2X0 U2486 ( .IN1(n1022), .IN2(n1632), .QN(g8766) );
  OA21X1 U2487 ( .IN1(g119), .IN2(n1633), .IN3(g109), .Q(g5918) );
  MUX21X1 U2488 ( .IN1(g1636), .IN2(g248), .S(g18), .Q(n1634) );
  INVX0 U2489 ( .INP(n1634), .ZN(n1842) );
  INVX0 U2490 ( .INP(g1462), .ZN(n1635) );
  OA221X1 U2491 ( .IN1(n1842), .IN2(n1635), .IN3(n1634), .IN4(g1462), .IN5(
        g109), .Q(g8045) );
  INVX0 U2492 ( .INP(g1806), .ZN(n1638) );
  OA221X1 U2493 ( .IN1(g1806), .IN2(n1639), .IN3(n1638), .IN4(n1637), .IN5(
        n1636), .Q(g8173) );
  MUX21X1 U2494 ( .IN1(g554), .IN2(g207), .S(g18), .Q(g6000) );
  INVX0 U2495 ( .INP(g158), .ZN(n1641) );
  INVX0 U2496 ( .INP(g6000), .ZN(n1640) );
  OA221X1 U2497 ( .IN1(g158), .IN2(g6000), .IN3(n1641), .IN4(n1640), .IN5(g109), .Q(g7843) );
  MUX21X1 U2498 ( .IN1(g572), .IN2(g243), .S(g18), .Q(g6042) );
  INVX0 U2499 ( .INP(g135), .ZN(n1643) );
  INVX0 U2500 ( .INP(g6042), .ZN(n1642) );
  OA221X1 U2501 ( .IN1(g135), .IN2(g6042), .IN3(n1643), .IN4(n1642), .IN5(g109), .Q(g8059) );
  INVX0 U2502 ( .INP(g1403), .ZN(n1644) );
  NAND2X0 U2503 ( .IN1(g18), .IN2(g207), .QN(n1652) );
  INVX0 U2504 ( .INP(n1652), .ZN(n1854) );
  MUX21X1 U2505 ( .IN1(n1644), .IN2(g1403), .S(n1854), .Q(n1645) );
  NOR2X0 U2506 ( .IN1(n1022), .IN2(n1645), .QN(g8767) );
  NOR2X0 U2507 ( .IN1(n1957), .IN2(n1646), .QN(n1647) );
  NOR2X0 U2508 ( .IN1(n1647), .IN2(g806), .QN(n1649) );
  NOR3X0 U2509 ( .IN1(n1649), .IN2(n1648), .IN3(n1817), .QN(g6126) );
  AND2X1 U2510 ( .IN1(n1669), .IN2(g631), .Q(g4891) );
  MUX21X1 U2511 ( .IN1(g546), .IN2(g186), .S(g18), .Q(g5996) );
  INVX0 U2512 ( .INP(g153), .ZN(n1683) );
  INVX0 U2513 ( .INP(g5996), .ZN(n1650) );
  OA221X1 U2514 ( .IN1(g153), .IN2(g5996), .IN3(n1683), .IN4(n1650), .IN5(g109), .Q(g8048) );
  INVX0 U2515 ( .INP(g1490), .ZN(n1651) );
  OA221X1 U2516 ( .IN1(n1652), .IN2(n1651), .IN3(n1854), .IN4(g1490), .IN5(
        g109), .Q(g8055) );
  INVX0 U2517 ( .INP(n1653), .ZN(n1654) );
  OAI22X1 U2518 ( .IN1(g105), .IN2(n1654), .IN3(n2023), .IN4(n1021), .QN(n1658) );
  NAND3X0 U2519 ( .IN1(g109), .IN2(g108), .IN3(g10722), .QN(n1656) );
  NAND3X0 U2520 ( .IN1(g109), .IN2(g865), .IN3(g10664), .QN(n1655) );
  NAND2X0 U2521 ( .IN1(n1656), .IN2(n1655), .QN(n1657) );
  NOR2X0 U2522 ( .IN1(n1658), .IN2(n1657), .QN(n2028) );
  AND2X1 U2523 ( .IN1(n2028), .IN2(g10515), .Q(g10583) );
  AND2X1 U2524 ( .IN1(g109), .IN2(g1362), .Q(g6820) );
  OA221X1 U2525 ( .IN1(n1661), .IN2(n1660), .IN3(n1659), .IN4(g1494), .IN5(
        g109), .Q(g8041) );
  AND2X1 U2526 ( .IN1(g109), .IN2(g248), .Q(g6840) );
  INVX0 U2527 ( .INP(n1662), .ZN(n1665) );
  OA221X1 U2528 ( .IN1(n1665), .IN2(g646), .IN3(n1665), .IN4(n1664), .IN5(
        n1663), .Q(g7134) );
  INVX0 U2529 ( .INP(n1666), .ZN(n1861) );
  MUX21X1 U2530 ( .IN1(n1667), .IN2(g1440), .S(n1861), .Q(n1668) );
  NOR2X0 U2531 ( .IN1(n1022), .IN2(n1668), .QN(g8772) );
  AND2X1 U2532 ( .IN1(n1669), .IN2(g635), .Q(g4893) );
  NAND2X0 U2533 ( .IN1(n1670), .IN2(n1945), .QN(n1671) );
  NOR4X0 U2534 ( .IN1(g617), .IN2(n1671), .IN3(n1940), .IN4(n1828), .QN(n1770)
         );
  NOR2X0 U2535 ( .IN1(n1770), .IN2(n1672), .QN(n1673) );
  MUX21X1 U2536 ( .IN1(g617), .IN2(n1941), .S(n1673), .Q(n1674) );
  NOR2X0 U2537 ( .IN1(n1606), .IN2(n1674), .QN(g8505) );
  INVX0 U2538 ( .INP(n1676), .ZN(n1678) );
  OA221X1 U2539 ( .IN1(g814), .IN2(n1678), .IN3(n1677), .IN4(n1676), .IN5(
        n1675), .Q(g7202) );
  MUX21X1 U2540 ( .IN1(g1811), .IN2(g201), .S(g18), .Q(n1815) );
  XOR3X1 U2541 ( .IN1(g1415), .IN2(g1515), .IN3(g1419), .Q(n1679) );
  XOR3X1 U2542 ( .IN1(n1815), .IN2(g1448), .IN3(n1679), .Q(n1680) );
  NOR2X0 U2543 ( .IN1(n1680), .IN2(n1022), .QN(g11514) );
  MUX21X1 U2544 ( .IN1(g1633), .IN2(g243), .S(g18), .Q(n1831) );
  INVX0 U2545 ( .INP(n1831), .ZN(n1682) );
  INVX0 U2546 ( .INP(g1466), .ZN(n1681) );
  OA221X1 U2547 ( .IN1(n1682), .IN2(n1681), .IN3(n1831), .IN4(g1466), .IN5(
        g109), .Q(g8051) );
  AND2X1 U2548 ( .IN1(g109), .IN2(g143), .Q(g6757) );
  NOR2X0 U2549 ( .IN1(g143), .IN2(n1022), .QN(n1685) );
  XNOR3X1 U2550 ( .IN1(g148), .IN2(g182), .IN3(n1683), .Q(n1684) );
  MUX21X1 U2551 ( .IN1(g6757), .IN2(n1685), .S(n1684), .Q(g6439) );
  NAND2X0 U2552 ( .IN1(g591), .IN2(g605), .QN(n1944) );
  INVX0 U2553 ( .INP(n1726), .ZN(n1725) );
  AO221X1 U2554 ( .IN1(g599), .IN2(g591), .IN3(n1778), .IN4(n1944), .IN5(n1725), .Q(n1686) );
  NAND2X0 U2555 ( .IN1(n1687), .IN2(n1686), .QN(n1688) );
  MUX21X1 U2556 ( .IN1(n1940), .IN2(g591), .S(n1688), .Q(n1689) );
  NOR2X0 U2557 ( .IN1(n1606), .IN2(n1689), .QN(g9110) );
  INVX0 U2558 ( .INP(g1478), .ZN(n1691) );
  OA221X1 U2559 ( .IN1(n1692), .IN2(n1691), .IN3(n1690), .IN4(g1478), .IN5(
        g109), .Q(g8043) );
  AND2X1 U2560 ( .IN1(g1848), .IN2(n1727), .Q(g4902) );
  NAND2X0 U2561 ( .IN1(n1694), .IN2(n1693), .QN(n1779) );
  INVX0 U2562 ( .INP(n1779), .ZN(n1695) );
  AO221X1 U2563 ( .IN1(g622), .IN2(n1991), .IN3(g622), .IN4(n1695), .IN5(n1705), .Q(g8820) );
  INVX0 U2564 ( .INP(g1436), .ZN(n1697) );
  MUX21X1 U2565 ( .IN1(g1436), .IN2(n1697), .S(n1696), .Q(n1698) );
  NOR2X0 U2566 ( .IN1(n1022), .IN2(n1698), .QN(g8775) );
  NOR2X0 U2567 ( .IN1(g1959), .IN2(n1008), .QN(n1700) );
  INVX0 U2568 ( .INP(n1700), .ZN(g4089) );
  OA21X1 U2569 ( .IN1(n2006), .IN2(n1881), .IN3(n1700), .Q(g5083) );
  NOR2X0 U2570 ( .IN1(g1696), .IN2(g4089), .QN(g5287) );
  MUX21X1 U2571 ( .IN1(g557), .IN2(g213), .S(g18), .Q(g6002) );
  INVX0 U2572 ( .INP(g162), .ZN(n1702) );
  INVX0 U2573 ( .INP(g6002), .ZN(n1701) );
  OA221X1 U2574 ( .IN1(g162), .IN2(g6002), .IN3(n1702), .IN4(n1701), .IN5(g109), .Q(g8060) );
  AND2X1 U2575 ( .IN1(g109), .IN2(g1411), .Q(g6244) );
  NOR3X0 U2576 ( .IN1(g591), .IN2(g599), .IN3(n1942), .QN(n1956) );
  OA221X1 U2577 ( .IN1(g591), .IN2(n1942), .IN3(n1940), .IN4(g605), .IN5(g599), 
        .Q(n1703) );
  OA21X1 U2578 ( .IN1(n1956), .IN2(n1703), .IN3(n1726), .Q(n1704) );
  NOR3X0 U2579 ( .IN1(n1961), .IN2(n1705), .IN3(n1704), .QN(n1706) );
  MUX21X1 U2580 ( .IN1(g605), .IN2(n1942), .S(n1706), .Q(n1707) );
  NOR2X0 U2581 ( .IN1(n1606), .IN2(n1707), .QN(g9150) );
  AND2X1 U2582 ( .IN1(g109), .IN2(g1504), .Q(g6215) );
  NAND4X0 U2583 ( .IN1(g1453), .IN2(g1494), .IN3(g1462), .IN4(g1508), .QN(
        n1713) );
  NAND3X0 U2584 ( .IN1(g1474), .IN2(g1478), .IN3(n1708), .QN(n1712) );
  INVX0 U2585 ( .INP(g1470), .ZN(n1719) );
  NOR4X0 U2586 ( .IN1(g1499), .IN2(g1482), .IN3(g1458), .IN4(n1719), .QN(n1709) );
  NAND4X0 U2587 ( .IN1(n1710), .IN2(n1709), .IN3(g1490), .IN4(g6215), .QN(
        n1711) );
  NOR4X0 U2588 ( .IN1(g1466), .IN2(n1713), .IN3(n1712), .IN4(n1711), .QN(n1714) );
  AO21X1 U2589 ( .IN1(g4), .IN2(g109), .IN3(n1714), .Q(g6656) );
  AND2X1 U2590 ( .IN1(g109), .IN2(g1371), .Q(g6824) );
  MUX21X1 U2591 ( .IN1(g575), .IN2(g248), .S(g18), .Q(g6045) );
  INVX0 U2592 ( .INP(g6045), .ZN(n1715) );
  OA221X1 U2593 ( .IN1(g139), .IN2(g6045), .IN3(n1716), .IN4(n1715), .IN5(g109), .Q(g8053) );
  OA221X1 U2594 ( .IN1(g1861), .IN2(g1845), .IN3(n1718), .IN4(n1717), .IN5(
        n1909), .Q(g6471) );
  MUX21X1 U2595 ( .IN1(g1630), .IN2(g237), .S(g18), .Q(n1966) );
  INVX0 U2596 ( .INP(n1966), .ZN(n1720) );
  OA221X1 U2597 ( .IN1(n1720), .IN2(n1719), .IN3(n1966), .IN4(g1470), .IN5(
        g109), .Q(g8039) );
  NOR2X0 U2598 ( .IN1(g758), .IN2(g762), .QN(n1723) );
  INVX0 U2599 ( .INP(n1721), .ZN(n1724) );
  NOR3X0 U2600 ( .IN1(n1723), .IN2(n1722), .IN3(n1724), .QN(g5529) );
  NOR2X0 U2601 ( .IN1(g758), .IN2(n1724), .QN(g4940) );
  OA221X1 U2602 ( .IN1(n1726), .IN2(g599), .IN3(n1725), .IN4(g605), .IN5(g18), 
        .Q(g9124) );
  AND2X1 U2603 ( .IN1(g109), .IN2(g231), .Q(g6822) );
  AND2X1 U2604 ( .IN1(g1853), .IN2(n1727), .Q(g4905) );
  OA221X1 U2605 ( .IN1(g466), .IN2(n1731), .IN3(n1730), .IN4(n1729), .IN5(
        n1728), .Q(g11376) );
  MUX21X1 U2606 ( .IN1(g995), .IN2(g1080), .S(n2007), .Q(g6895) );
  AO22X1 U2607 ( .IN1(n1289), .IN2(g1235), .IN3(g1240), .IN4(n2010), .Q(g7297)
         );
  MUX21X1 U2608 ( .IN1(g1621), .IN2(n1854), .S(n2007), .Q(g8771) );
  OA21X1 U2609 ( .IN1(g1840), .IN2(n1795), .IN3(n1733), .Q(n1998) );
  NOR2X0 U2610 ( .IN1(n1749), .IN2(n1998), .QN(n1997) );
  NAND2X0 U2611 ( .IN1(n1735), .IN2(n1734), .QN(n1736) );
  AO22X1 U2612 ( .IN1(n1998), .IN2(g1950), .IN3(n1997), .IN4(n1736), .Q(n1737)
         );
  MUX21X1 U2613 ( .IN1(g1945), .IN2(n1738), .S(n1737), .Q(n1742) );
  NOR2X0 U2614 ( .IN1(n2002), .IN2(n1740), .QN(n1741) );
  AO21X1 U2615 ( .IN1(n2002), .IN2(n1742), .IN3(n1741), .Q(g8945) );
  AO22X1 U2616 ( .IN1(g727), .IN2(n2004), .IN3(g736), .IN4(n2003), .Q(g8435)
         );
  MUX21X1 U2617 ( .IN1(g135), .IN2(g293), .S(n2005), .Q(g6911) );
  MUX21X1 U2618 ( .IN1(g991), .IN2(g1083), .S(n2007), .Q(g6898) );
  MUX21X1 U2619 ( .IN1(g178), .IN2(g266), .S(n2005), .Q(g6900) );
  MUX21X1 U2620 ( .IN1(g1092), .IN2(g360), .S(n2006), .Q(g6088) );
  MUX21X1 U2621 ( .IN1(g166), .IN2(g299), .S(n2005), .Q(g6923) );
  OR2X1 U2622 ( .IN1(n1743), .IN2(n1022), .Q(n1745) );
  NAND2X0 U2623 ( .IN1(n1745), .IN2(n1744), .QN(n1746) );
  MUX21X1 U2624 ( .IN1(g947), .IN2(g833), .S(n1934), .Q(g11300) );
  AO21X1 U2625 ( .IN1(g1681), .IN2(n1971), .IN3(n1748), .Q(g10864) );
  MUX21X1 U2626 ( .IN1(g1098), .IN2(g366), .S(n2006), .Q(g6096) );
  MUX21X1 U2627 ( .IN1(g968), .IN2(g861), .S(n1934), .Q(g11314) );
  INVX0 U2628 ( .INP(n1998), .ZN(n1757) );
  NAND2X0 U2629 ( .IN1(n1749), .IN2(n1757), .QN(n1929) );
  OA21X1 U2630 ( .IN1(g1878), .IN2(n1757), .IN3(n1929), .Q(n1750) );
  MUX21X1 U2631 ( .IN1(g1872), .IN2(n1489), .S(n1750), .Q(n1751) );
  AO21X1 U2632 ( .IN1(n2002), .IN2(n1751), .IN3(n1741), .Q(g8921) );
  MUX21X1 U2633 ( .IN1(g1436), .IN2(g1598), .S(n1992), .Q(g6481) );
  MUX21X1 U2634 ( .IN1(n1752), .IN2(g366), .S(n2008), .Q(g11487) );
  INVX0 U2635 ( .INP(g1927), .ZN(n1761) );
  INVX0 U2636 ( .INP(g1932), .ZN(n1758) );
  NAND2X0 U2637 ( .IN1(n1753), .IN2(n1757), .QN(n1845) );
  OR2X1 U2638 ( .IN1(n1998), .IN2(n1754), .Q(n1844) );
  OAI222X1 U2639 ( .IN1(n1758), .IN2(n1757), .IN3(n1845), .IN4(n1756), .IN5(
        n1844), .IN6(n1755), .QN(n1759) );
  NAND2X0 U2640 ( .IN1(n1929), .IN2(n1759), .QN(n1760) );
  MUX21X1 U2641 ( .IN1(n1761), .IN2(g1927), .S(n1760), .Q(n1762) );
  AO21X1 U2642 ( .IN1(n2002), .IN2(n1762), .IN3(n1741), .Q(g8941) );
  OAI21X1 U2643 ( .IN1(n1288), .IN2(n1765), .IN3(n1764), .QN(n1766) );
  AO22X1 U2644 ( .IN1(n1766), .IN2(n1289), .IN3(g1275), .IN4(n1028), .Q(g11443) );
  AO22X1 U2645 ( .IN1(g700), .IN2(n2003), .IN3(g691), .IN4(n2004), .Q(g8431)
         );
  AO221X1 U2646 ( .IN1(g1766), .IN2(n1768), .IN3(n1767), .IN4(n1881), .IN5(
        g1713), .Q(g7133) );
  AO22X1 U2647 ( .IN1(g1923), .IN2(n1915), .IN3(g1932), .IN4(n1916), .Q(g8286)
         );
  AO22X1 U2648 ( .IN1(n1289), .IN2(g1270), .IN3(g1304), .IN4(n2010), .Q(g7290)
         );
  MUX21X1 U2649 ( .IN1(g1083), .IN2(g351), .S(n2006), .Q(g6068) );
  MUX21X1 U2650 ( .IN1(g1415), .IN2(g1567), .S(n1992), .Q(g6468) );
  MUX21X1 U2651 ( .IN1(n1769), .IN2(g339), .S(n2008), .Q(g11478) );
  AO22X1 U2652 ( .IN1(g1932), .IN2(n1915), .IN3(g1941), .IN4(n1916), .Q(g8287)
         );
  MUX21X1 U2653 ( .IN1(g1428), .IN2(g1589), .S(n1992), .Q(g6524) );
  MUX21X1 U2654 ( .IN1(g1032), .IN2(g1077), .S(n2007), .Q(g7257) );
  AO22X1 U2655 ( .IN1(n1289), .IN2(g1255), .IN3(g1260), .IN4(n2010), .Q(g7301)
         );
  MUX21X1 U2656 ( .IN1(g496), .IN2(g501), .S(n1968), .Q(g11334) );
  NOR2X0 U2657 ( .IN1(n1771), .IN2(n1770), .QN(n1871) );
  NAND2X0 U2658 ( .IN1(n1773), .IN2(n1772), .QN(n1775) );
  NOR2X0 U2659 ( .IN1(n1986), .IN2(n1774), .QN(n1937) );
  INVX0 U2660 ( .INP(n1937), .ZN(n1985) );
  OA221X1 U2661 ( .IN1(n1871), .IN2(g727), .IN3(n1986), .IN4(n1775), .IN5(
        n1985), .Q(n1776) );
  MUX21X1 U2662 ( .IN1(g722), .IN2(n1777), .S(n1776), .Q(n1780) );
  NOR2X0 U2663 ( .IN1(g605), .IN2(n1778), .QN(n1951) );
  NOR4X0 U2664 ( .IN1(n1991), .IN2(n1951), .IN3(n1956), .IN4(n1779), .QN(n1989) );
  AO21X1 U2665 ( .IN1(n1991), .IN2(n1780), .IN3(n1989), .Q(g8923) );
  INVX0 U2666 ( .INP(g1718), .ZN(n1967) );
  NAND2X0 U2667 ( .IN1(n1781), .IN2(n1967), .QN(n1782) );
  NOR2X0 U2668 ( .IN1(n1782), .IN2(n1971), .QN(n1841) );
  AO21X1 U2669 ( .IN1(g566), .IN2(n1971), .IN3(n1841), .Q(g10799) );
  AO21X1 U2670 ( .IN1(g563), .IN2(n1971), .IN3(n1783), .Q(g10798) );
  MUX21X1 U2671 ( .IN1(n1489), .IN2(g1872), .S(n1784), .Q(n1785) );
  AO22X1 U2672 ( .IN1(n1998), .IN2(g1887), .IN3(n1997), .IN4(n1785), .Q(n1786)
         );
  MUX21X1 U2673 ( .IN1(g1882), .IN2(n1490), .S(n1786), .Q(n1787) );
  AO21X1 U2674 ( .IN1(n2002), .IN2(n1787), .IN3(n1741), .Q(g8943) );
  INVX0 U2675 ( .INP(g1690), .ZN(n2013) );
  NOR2X0 U2676 ( .IN1(g10719), .IN2(n2013), .QN(n1803) );
  NOR2X0 U2677 ( .IN1(g1690), .IN2(g1806), .QN(n1802) );
  NOR2X0 U2678 ( .IN1(g1822), .IN2(g1834), .QN(n1789) );
  NAND2X0 U2679 ( .IN1(n1789), .IN2(n1788), .QN(n1796) );
  NOR2X0 U2680 ( .IN1(g1834), .IN2(n1790), .QN(n1792) );
  MUX21X1 U2681 ( .IN1(n1792), .IN2(n1791), .S(g1857), .Q(n1794) );
  NOR2X0 U2682 ( .IN1(n1022), .IN2(g10724), .QN(n1912) );
  NAND2X0 U2683 ( .IN1(n1794), .IN2(n1912), .QN(n1793) );
  OA221X1 U2684 ( .IN1(n1796), .IN2(n1795), .IN3(n1794), .IN4(n1912), .IN5(
        n1793), .Q(n1797) );
  NAND2X0 U2685 ( .IN1(g4904), .IN2(n1797), .QN(n1800) );
  INVX0 U2686 ( .INP(n1798), .ZN(n1799) );
  AO21X1 U2687 ( .IN1(g1854), .IN2(n1800), .IN3(n1799), .Q(n1801) );
  AO222X1 U2688 ( .IN1(n1804), .IN2(n1803), .IN3(n1804), .IN4(n1802), .IN5(
        n1903), .IN6(n1801), .Q(g11293) );
  MUX21X1 U2689 ( .IN1(g391), .IN2(g396), .S(n1968), .Q(g11265) );
  INVX0 U2690 ( .INP(g695), .ZN(n1863) );
  INVX0 U2691 ( .INP(g658), .ZN(n1857) );
  NAND2X0 U2692 ( .IN1(n1871), .IN2(n1806), .QN(n1983) );
  INVX0 U2693 ( .INP(g677), .ZN(n1808) );
  INVX0 U2694 ( .INP(g668), .ZN(n1807) );
  NAND2X0 U2695 ( .IN1(n1808), .IN2(n1807), .QN(n1809) );
  NOR2X0 U2696 ( .IN1(n1983), .IN2(n1809), .QN(n1883) );
  NAND3X0 U2697 ( .IN1(g658), .IN2(n1871), .IN3(n1810), .QN(n1984) );
  NOR2X0 U2698 ( .IN1(n1811), .IN2(n1984), .QN(n1918) );
  MUX21X1 U2699 ( .IN1(n1883), .IN2(n1918), .S(g686), .Q(n1812) );
  OA221X1 U2700 ( .IN1(n1812), .IN2(g700), .IN3(n1812), .IN4(n1986), .IN5(
        n1985), .Q(n1813) );
  MUX21X1 U2701 ( .IN1(g695), .IN2(n1863), .S(n1813), .Q(n1814) );
  AO21X1 U2702 ( .IN1(n1991), .IN2(n1814), .IN3(n1989), .Q(g8887) );
  MUX21X1 U2703 ( .IN1(g1407), .IN2(g1586), .S(n1992), .Q(g6514) );
  AO22X1 U2704 ( .IN1(g709), .IN2(n2004), .IN3(g718), .IN4(n2003), .Q(g8433)
         );
  MUX21X1 U2705 ( .IN1(g1618), .IN2(n1815), .S(n2007), .Q(g11579) );
  MUX21X1 U2706 ( .IN1(n1816), .IN2(g1724), .S(n1913), .Q(g10771) );
  MUX21X1 U2707 ( .IN1(g1504), .IN2(g1528), .S(n1992), .Q(g6522) );
  AO221X1 U2708 ( .IN1(n1957), .IN2(g798), .IN3(n1957), .IN4(g794), .IN5(n1817), .Q(g6243) );
  MUX21X1 U2709 ( .IN1(g1458), .IN2(g1561), .S(n1992), .Q(g6542) );
  AO22X1 U2710 ( .IN1(n1289), .IN2(g1265), .IN3(g1270), .IN4(n2010), .Q(g7303)
         );
  MUX21X1 U2711 ( .IN1(g1003), .IN2(g1086), .S(n2007), .Q(g6902) );
  MUX21X1 U2712 ( .IN1(g1470), .IN2(g1552), .S(n1992), .Q(g6529) );
  MUX21X1 U2713 ( .IN1(g386), .IN2(g391), .S(n1964), .Q(g11264) );
  NAND2X0 U2714 ( .IN1(n1818), .IN2(n1967), .QN(n1819) );
  NOR2X0 U2715 ( .IN1(n1819), .IN2(n1971), .QN(n1926) );
  AO21X1 U2716 ( .IN1(g557), .IN2(n1971), .IN3(n1926), .Q(g10795) );
  MUX21X1 U2717 ( .IN1(g1791), .IN2(g1324), .S(n1965), .Q(g11607) );
  MUX21X1 U2718 ( .IN1(g1657), .IN2(g1675), .S(g1690), .Q(g3414) );
  AO22X1 U2719 ( .IN1(n1289), .IN2(g1292), .IN3(g1284), .IN4(n2010), .Q(g7294)
         );
  NOR2X0 U2720 ( .IN1(g1900), .IN2(n1844), .QN(n1928) );
  NOR2X0 U2721 ( .IN1(n1848), .IN2(n1845), .QN(n1927) );
  NOR2X0 U2722 ( .IN1(n1928), .IN2(n1927), .QN(n1821) );
  NAND2X0 U2723 ( .IN1(n1998), .IN2(g1914), .QN(n1820) );
  NAND2X0 U2724 ( .IN1(n1821), .IN2(n1820), .QN(n1822) );
  NAND2X0 U2725 ( .IN1(n1929), .IN2(n1822), .QN(n1823) );
  MUX21X1 U2726 ( .IN1(n1824), .IN2(g1909), .S(n1823), .Q(n1825) );
  AO21X1 U2727 ( .IN1(n2002), .IN2(n1825), .IN3(n1741), .Q(g8939) );
  MUX21X1 U2728 ( .IN1(g538), .IN2(g534), .S(n1964), .Q(g11327) );
  MUX21X1 U2729 ( .IN1(g1786), .IN2(g1321), .S(n1965), .Q(g11606) );
  MUX21X1 U2730 ( .IN1(g950), .IN2(g837), .S(n1934), .Q(g11303) );
  MUX21X1 U2731 ( .IN1(g1424), .IN2(g1583), .S(n1992), .Q(g6506) );
  NOR2X0 U2732 ( .IN1(n1828), .IN2(g639), .QN(n1827) );
  AO221X1 U2733 ( .IN1(g639), .IN2(n1828), .IN3(n1827), .IN4(n1826), .IN5(
        n1961), .Q(g7626) );
  MUX21X1 U2734 ( .IN1(n1829), .IN2(g1721), .S(n1913), .Q(g10770) );
  MUX21X1 U2735 ( .IN1(n1830), .IN2(g354), .S(n2008), .Q(g11483) );
  MUX21X1 U2736 ( .IN1(g1482), .IN2(g1543), .S(n1992), .Q(g6545) );
  OR2X1 U2737 ( .IN1(g1718), .IN2(n1831), .Q(n1839) );
  MUX21X1 U2738 ( .IN1(n1839), .IN2(g1657), .S(n1978), .Q(g10767) );
  MUX21X1 U2739 ( .IN1(g542), .IN2(g538), .S(n1968), .Q(g11326) );
  MUX21X1 U2740 ( .IN1(g1027), .IN2(n1832), .S(g999), .Q(n1834) );
  XNOR3X1 U2741 ( .IN1(g1023), .IN2(g1015), .IN3(g1007), .Q(n1833) );
  XNOR3X1 U2742 ( .IN1(g1003), .IN2(n1834), .IN3(n1833), .Q(n1835) );
  XNOR3X1 U2743 ( .IN1(g1019), .IN2(g1011), .IN3(n1835), .Q(n1836) );
  XNOR3X1 U2744 ( .IN1(g991), .IN2(g995), .IN3(n1836), .Q(n1837) );
  AO222X1 U2745 ( .IN1(n2007), .IN2(n1838), .IN3(n2007), .IN4(n1837), .IN5(
        g105), .IN6(n1971), .Q(g10898) );
  MUX21X1 U2746 ( .IN1(g1444), .IN2(g1604), .S(n1992), .Q(g6507) );
  MUX21X1 U2747 ( .IN1(g572), .IN2(n1839), .S(n2007), .Q(g10718) );
  AO22X1 U2748 ( .IN1(n1289), .IN2(g1300), .IN3(g1296), .IN4(n2010), .Q(g7292)
         );
  OR2X1 U2749 ( .IN1(g1718), .IN2(n1840), .Q(n1859) );
  MUX21X1 U2750 ( .IN1(n1859), .IN2(g1663), .S(n1978), .Q(g10861) );
  AO21X1 U2751 ( .IN1(g1687), .IN2(n1971), .IN3(n1841), .Q(g10776) );
  NAND2X0 U2752 ( .IN1(n1967), .IN2(n1842), .QN(n1875) );
  MUX21X1 U2753 ( .IN1(n1875), .IN2(g1660), .S(n1978), .Q(g10859) );
  AO22X1 U2754 ( .IN1(n1289), .IN2(g1245), .IN3(g1250), .IN4(n2010), .Q(g7299)
         );
  AO21X1 U2755 ( .IN1(g1672), .IN2(n1971), .IN3(n1843), .Q(g10858) );
  MUX21X1 U2756 ( .IN1(g1023), .IN2(g1071), .S(n2007), .Q(g7244) );
  MUX21X1 U2757 ( .IN1(g1660), .IN2(g1678), .S(g1690), .Q(g3425) );
  MUX21X1 U2758 ( .IN1(g999), .IN2(g1089), .S(n2007), .Q(g6908) );
  NAND2X0 U2759 ( .IN1(n1845), .IN2(n1844), .QN(n1846) );
  OA221X1 U2760 ( .IN1(n1846), .IN2(n1998), .IN3(n1846), .IN4(g1905), .IN5(
        n1929), .Q(n1847) );
  MUX21X1 U2761 ( .IN1(g1900), .IN2(n1848), .S(n1847), .Q(n1849) );
  AO21X1 U2762 ( .IN1(n2002), .IN2(n1849), .IN3(n1741), .Q(g8938) );
  MUX21X1 U2763 ( .IN1(g1071), .IN2(g339), .S(n2006), .Q(g5910) );
  MUX21X1 U2764 ( .IN1(n1850), .IN2(g351), .S(n2008), .Q(g11482) );
  MUX21X1 U2765 ( .IN1(g1713), .IN2(g1710), .S(n2007), .Q(g5396) );
  AO22X1 U2766 ( .IN1(n1289), .IN2(g1284), .IN3(g1280), .IN4(n1028), .Q(g7295)
         );
  AO22X1 U2767 ( .IN1(g1914), .IN2(n1916), .IN3(g1905), .IN4(n1915), .Q(g8284)
         );
  MUX21X1 U2768 ( .IN1(g127), .IN2(g287), .S(n2005), .Q(g6901) );
  NAND2X0 U2769 ( .IN1(g1878), .IN2(n1851), .QN(n1852) );
  NAND3X0 U2770 ( .IN1(n1903), .IN2(n1853), .IN3(n1852), .QN(g8559) );
  NOR2X0 U2771 ( .IN1(g1718), .IN2(n1854), .QN(n1855) );
  NOR2X0 U2772 ( .IN1(n1971), .IN2(n1855), .QN(n1970) );
  AO21X1 U2773 ( .IN1(g1675), .IN2(n1971), .IN3(n1970), .Q(g10860) );
  OA21X1 U2774 ( .IN1(n1871), .IN2(g664), .IN3(n1985), .Q(n1856) );
  MUX21X1 U2775 ( .IN1(g658), .IN2(n1857), .S(n1856), .Q(n1858) );
  AO21X1 U2776 ( .IN1(n1991), .IN2(n1858), .IN3(n1989), .Q(g8973) );
  MUX21X1 U2777 ( .IN1(g1411), .IN2(g1580), .S(n1992), .Q(g6500) );
  MUX21X1 U2778 ( .IN1(g549), .IN2(n1859), .S(n2007), .Q(g10855) );
  MUX21X1 U2779 ( .IN1(g1771), .IN2(g1311), .S(n1965), .Q(g11603) );
  OR2X1 U2780 ( .IN1(g627), .IN2(n1005), .Q(g6672) );
  MUX21X1 U2781 ( .IN1(g1474), .IN2(g1549), .S(n1992), .Q(g6523) );
  INVX0 U2782 ( .INP(n1876), .ZN(n1860) );
  MUX21X1 U2783 ( .IN1(n1860), .IN2(g1730), .S(n1913), .Q(g10707) );
  AO22X1 U2784 ( .IN1(n1289), .IN2(g1240), .IN3(g1245), .IN4(n1028), .Q(g7298)
         );
  MUX21X1 U2785 ( .IN1(g1478), .IN2(g1546), .S(n1992), .Q(g6551) );
  MUX21X1 U2786 ( .IN1(g1074), .IN2(g342), .S(n2006), .Q(g6099) );
  AO22X1 U2787 ( .IN1(g1887), .IN2(n1915), .IN3(g1896), .IN4(n1916), .Q(g8282)
         );
  MUX21X1 U2788 ( .IN1(g1466), .IN2(g1555), .S(n1992), .Q(g6534) );
  MUX21X1 U2789 ( .IN1(g1630), .IN2(n1861), .S(n2007), .Q(g8776) );
  MUX21X1 U2790 ( .IN1(g1508), .IN2(g1524), .S(n1992), .Q(g6513) );
  MUX21X1 U2791 ( .IN1(g139), .IN2(g296), .S(n2005), .Q(g6916) );
  MUX21X1 U2792 ( .IN1(g1633), .IN2(n1862), .S(n2007), .Q(g8777) );
  AO22X1 U2793 ( .IN1(n1289), .IN2(g1304), .IN3(g1300), .IN4(n1028), .Q(g7291)
         );
  MUX21X1 U2794 ( .IN1(g525), .IN2(g521), .S(n1964), .Q(g11330) );
  MUX21X1 U2795 ( .IN1(g1077), .IN2(g345), .S(n2006), .Q(g5914) );
  MUX21X1 U2796 ( .IN1(g452), .IN2(g448), .S(n1964), .Q(g11258) );
  MUX21X1 U2797 ( .IN1(g1068), .IN2(g336), .S(n2006), .Q(g6054) );
  MUX21X1 U2798 ( .IN1(g1766), .IN2(g1308), .S(n1965), .Q(g11602) );
  MUX21X1 U2799 ( .IN1(g511), .IN2(g516), .S(n1964), .Q(g11337) );
  INVX0 U2800 ( .INP(g686), .ZN(n1888) );
  AND3X1 U2801 ( .IN1(n1883), .IN2(n1888), .IN3(n1863), .Q(n1920) );
  NOR2X0 U2802 ( .IN1(n1888), .IN2(n1863), .QN(n1864) );
  AO22X1 U2803 ( .IN1(n1864), .IN2(n1918), .IN3(g709), .IN4(n1986), .Q(n1865)
         );
  OA21X1 U2804 ( .IN1(n1920), .IN2(n1865), .IN3(n1985), .Q(n1866) );
  MUX21X1 U2805 ( .IN1(g704), .IN2(n1921), .S(n1866), .Q(n1867) );
  AO21X1 U2806 ( .IN1(n1991), .IN2(n1867), .IN3(n1989), .Q(g8889) );
  AO22X1 U2807 ( .IN1(g1923), .IN2(n1916), .IN3(g1914), .IN4(n1915), .Q(g8285)
         );
  MUX21X1 U2808 ( .IN1(g506), .IN2(g511), .S(n1968), .Q(g11336) );
  OR2X1 U2809 ( .IN1(n1869), .IN2(n1868), .Q(n1870) );
  OA221X1 U2810 ( .IN1(n1871), .IN2(g736), .IN3(n1986), .IN4(n1870), .IN5(
        n1985), .Q(n1872) );
  MUX21X1 U2811 ( .IN1(g731), .IN2(n1873), .S(n1872), .Q(n1874) );
  AO21X1 U2812 ( .IN1(n1991), .IN2(n1874), .IN3(n1989), .Q(g8926) );
  AO22X1 U2813 ( .IN1(n1289), .IN2(g1296), .IN3(g1292), .IN4(n1028), .Q(g7293)
         );
  MUX21X1 U2814 ( .IN1(g575), .IN2(n1875), .S(n2007), .Q(g10800) );
  MUX21X1 U2815 ( .IN1(g959), .IN2(g849), .S(n1934), .Q(g11308) );
  NAND3X0 U2816 ( .IN1(n1880), .IN2(n1879), .IN3(n1878), .QN(n1882) );
  MUX21X1 U2817 ( .IN1(g1811), .IN2(n1882), .S(n1881), .Q(g10936) );
  MUX21X1 U2818 ( .IN1(g1403), .IN2(g1592), .S(n1992), .Q(g6470) );
  MUX21X1 U2819 ( .IN1(g182), .IN2(g263), .S(n2005), .Q(g6897) );
  NOR2X0 U2820 ( .IN1(n1883), .IN2(n1918), .QN(n1885) );
  NAND2X0 U2821 ( .IN1(g691), .IN2(n1986), .QN(n1884) );
  NAND2X0 U2822 ( .IN1(n1885), .IN2(n1884), .QN(n1886) );
  NAND2X0 U2823 ( .IN1(n1985), .IN2(n1886), .QN(n1887) );
  MUX21X1 U2824 ( .IN1(n1888), .IN2(g686), .S(n1887), .Q(n1889) );
  AO21X1 U2825 ( .IN1(n1991), .IN2(n1889), .IN3(n1989), .Q(g8885) );
  MUX21X1 U2826 ( .IN1(n1890), .IN2(g342), .S(n2008), .Q(g11488) );
  AO22X1 U2827 ( .IN1(g1950), .IN2(n1916), .IN3(g1941), .IN4(n1915), .Q(g8288)
         );
  MUX21X1 U2828 ( .IN1(g1806), .IN2(g1333), .S(n1965), .Q(g11610) );
  MUX21X1 U2829 ( .IN1(g416), .IN2(g421), .S(n1968), .Q(g11270) );
  MUX21X1 U2830 ( .IN1(g1080), .IN2(g348), .S(n2006), .Q(g6059) );
  NOR2X0 U2831 ( .IN1(n1892), .IN2(n1891), .QN(n1907) );
  NAND2X0 U2832 ( .IN1(g10724), .IN2(n2029), .QN(n1893) );
  NAND2X0 U2833 ( .IN1(n1893), .IN2(g1690), .QN(n1895) );
  AO21X1 U2834 ( .IN1(g1786), .IN2(g1791), .IN3(g1690), .Q(n1894) );
  AND2X1 U2835 ( .IN1(n1895), .IN2(n1894), .Q(n1902) );
  AO21X1 U2836 ( .IN1(g1766), .IN2(g1771), .IN3(g1690), .Q(n1896) );
  OA221X1 U2837 ( .IN1(n2013), .IN2(g10719), .IN3(n2013), .IN4(g10720), .IN5(
        n1896), .Q(n1900) );
  NOR2X0 U2838 ( .IN1(n1900), .IN2(n1897), .QN(n1898) );
  NOR2X0 U2839 ( .IN1(n1898), .IN2(n2013), .QN(n1899) );
  OA221X1 U2840 ( .IN1(n1902), .IN2(g10664), .IN3(n1902), .IN4(g10663), .IN5(
        n1899), .Q(n1905) );
  OA221X1 U2841 ( .IN1(n1900), .IN2(g1776), .IN3(n1900), .IN4(g1781), .IN5(
        n2013), .Q(n1901) );
  OA221X1 U2842 ( .IN1(n1902), .IN2(g1796), .IN3(n1902), .IN4(g1801), .IN5(
        n1901), .Q(n1904) );
  NOR3X0 U2843 ( .IN1(n1905), .IN2(n1904), .IN3(n1903), .QN(n1906) );
  AO221X1 U2844 ( .IN1(g1857), .IN2(n1909), .IN3(n1908), .IN4(n1907), .IN5(
        n1906), .Q(g11294) );
  OA21X1 U2845 ( .IN1(n2007), .IN2(g1718), .IN3(n1910), .Q(g5404) );
  MUX21X1 U2846 ( .IN1(g1718), .IN2(g1666), .S(n1978), .Q(g10863) );
  AO22X1 U2847 ( .IN1(g682), .IN2(n2003), .IN3(g673), .IN4(n2004), .Q(g8429)
         );
  AO22X1 U2848 ( .IN1(g1878), .IN2(n1915), .IN3(g1887), .IN4(n1916), .Q(g8281)
         );
  MUX21X1 U2849 ( .IN1(g153), .IN2(g272), .S(n2005), .Q(g6910) );
  MUX21X1 U2850 ( .IN1(g953), .IN2(g841), .S(n1934), .Q(g11305) );
  MUX21X1 U2851 ( .IN1(g1462), .IN2(g1558), .S(n1992), .Q(g6538) );
  MUX21X1 U2852 ( .IN1(g1095), .IN2(g363), .S(n2006), .Q(g6093) );
  MUX21X1 U2853 ( .IN1(n1911), .IN2(g360), .S(n2008), .Q(g11485) );
  MUX21X1 U2854 ( .IN1(g1666), .IN2(g1684), .S(g1690), .Q(g3435) );
  INVX0 U2855 ( .INP(n1912), .ZN(n1914) );
  MUX21X1 U2856 ( .IN1(n1914), .IN2(g1733), .S(n1913), .Q(g10711) );
  AO22X1 U2857 ( .IN1(g1905), .IN2(n1916), .IN3(g1896), .IN4(n1915), .Q(g8283)
         );
  INVX0 U2858 ( .INP(g713), .ZN(n1924) );
  INVX0 U2859 ( .INP(n1917), .ZN(n1919) );
  AO222X1 U2860 ( .IN1(n1921), .IN2(n1920), .IN3(n1986), .IN4(g718), .IN5(
        n1919), .IN6(n1918), .Q(n1922) );
  NAND2X0 U2861 ( .IN1(n1985), .IN2(n1922), .QN(n1923) );
  MUX21X1 U2862 ( .IN1(n1924), .IN2(g713), .S(n1923), .Q(n1925) );
  AO21X1 U2863 ( .IN1(n1991), .IN2(n1925), .IN3(n1989), .Q(g8920) );
  AO21X1 U2864 ( .IN1(g1678), .IN2(n1971), .IN3(n1926), .Q(g10862) );
  MUX21X1 U2865 ( .IN1(g491), .IN2(g496), .S(n1968), .Q(g11333) );
  MUX21X1 U2866 ( .IN1(g1089), .IN2(g357), .S(n2006), .Q(g6080) );
  MUX21X1 U2867 ( .IN1(g1419), .IN2(g1577), .S(n1992), .Q(g6480) );
  MUX21X1 U2868 ( .IN1(g1801), .IN2(g1330), .S(n1965), .Q(g11609) );
  MUX21X1 U2869 ( .IN1(n1928), .IN2(n1927), .S(g1909), .Q(n1930) );
  OA221X1 U2870 ( .IN1(n1930), .IN2(n1998), .IN3(n1930), .IN4(g1923), .IN5(
        n1929), .Q(n1931) );
  MUX21X1 U2871 ( .IN1(g1918), .IN2(n1932), .S(n1931), .Q(n1933) );
  AO21X1 U2872 ( .IN1(n2002), .IN2(n1933), .IN3(n1741), .Q(g8940) );
  MUX21X1 U2873 ( .IN1(n1019), .IN2(g857), .S(n1934), .Q(g11312) );
  AO22X1 U2874 ( .IN1(g673), .IN2(n2003), .IN3(g664), .IN4(n2004), .Q(g8428)
         );
  AO22X1 U2875 ( .IN1(g691), .IN2(n2003), .IN3(g682), .IN4(n2004), .Q(g8430)
         );
  MUX21X1 U2876 ( .IN1(g1019), .IN2(g1098), .S(n2007), .Q(g6924) );
  NAND2X0 U2877 ( .IN1(g682), .IN2(n1986), .QN(n1935) );
  OA221X1 U2878 ( .IN1(g668), .IN2(n1983), .IN3(n1807), .IN4(n1984), .IN5(
        n1935), .Q(n1936) );
  NOR2X0 U2879 ( .IN1(n1937), .IN2(n1936), .QN(n1938) );
  MUX21X1 U2880 ( .IN1(g677), .IN2(n1808), .S(n1938), .Q(n1939) );
  AO21X1 U2881 ( .IN1(n1991), .IN2(n1939), .IN3(n1989), .Q(g8883) );
  MUX21X1 U2882 ( .IN1(g530), .IN2(g525), .S(n1964), .Q(g11329) );
  MUX21X1 U2883 ( .IN1(g534), .IN2(g530), .S(n1964), .Q(g11328) );
  AO22X1 U2884 ( .IN1(n1289), .IN2(g1250), .IN3(g1255), .IN4(n1028), .Q(g7300)
         );
  MUX21X1 U2885 ( .IN1(g1494), .IN2(g1534), .S(n1992), .Q(g6533) );
  MUX21X1 U2886 ( .IN1(g1663), .IN2(g1681), .S(g1690), .Q(g3431) );
  INVX0 U2887 ( .INP(g622), .ZN(n1955) );
  NAND2X0 U2888 ( .IN1(g599), .IN2(n1940), .QN(n1946) );
  NAND2X0 U2889 ( .IN1(n1942), .IN2(n1941), .QN(n1943) );
  NAND4X0 U2890 ( .IN1(n1945), .IN2(n1946), .IN3(n1944), .IN4(n1943), .QN(
        n1952) );
  NAND2X0 U2891 ( .IN1(g622), .IN2(g255), .QN(n1950) );
  AND2X1 U2892 ( .IN1(n1945), .IN2(n1944), .Q(n1947) );
  MUX21X1 U2893 ( .IN1(n1947), .IN2(n1946), .S(g639), .Q(n1949) );
  NAND2X0 U2894 ( .IN1(n1950), .IN2(n1949), .QN(n1948) );
  OA221X1 U2895 ( .IN1(n1952), .IN2(n1951), .IN3(n1950), .IN4(n1949), .IN5(
        n1948), .Q(n1953) );
  NAND2X0 U2896 ( .IN1(g4892), .IN2(n1953), .QN(n1954) );
  AO22X1 U2897 ( .IN1(n1956), .IN2(n1955), .IN3(g636), .IN4(n1954), .Q(n1963)
         );
  NAND2X0 U2898 ( .IN1(n1958), .IN2(n1957), .QN(n1960) );
  AO22X1 U2899 ( .IN1(g810), .IN2(g814), .IN3(g818), .IN4(g822), .Q(n1959) );
  NAND3X0 U2900 ( .IN1(n1960), .IN2(n1959), .IN3(g826), .QN(n1962) );
  MUX21X1 U2901 ( .IN1(n1963), .IN2(n1962), .S(n1961), .Q(g8631) );
  MUX21X1 U2902 ( .IN1(g162), .IN2(g278), .S(n2005), .Q(g6922) );
  MUX21X1 U2903 ( .IN1(g426), .IN2(g386), .S(n1964), .Q(g11263) );
  MUX21X1 U2904 ( .IN1(g1432), .IN2(g1595), .S(n1992), .Q(g6479) );
  MUX21X1 U2905 ( .IN1(g1440), .IN2(g1601), .S(n1992), .Q(g6501) );
  MUX21X1 U2906 ( .IN1(g1654), .IN2(g1672), .S(g1690), .Q(g3399) );
  MUX21X1 U2907 ( .IN1(g1781), .IN2(g1318), .S(n1965), .Q(g11605) );
  AND2X1 U2908 ( .IN1(n1967), .IN2(n1966), .Q(n1979) );
  MUX21X1 U2909 ( .IN1(g569), .IN2(n1979), .S(n2007), .Q(g10717) );
  MUX21X1 U2910 ( .IN1(g1011), .IN2(g1092), .S(n2007), .Q(g6912) );
  MUX21X1 U2911 ( .IN1(g143), .IN2(g302), .S(n2005), .Q(g6929) );
  MUX21X1 U2912 ( .IN1(g476), .IN2(g542), .S(n1968), .Q(g11325) );
  MUX21X1 U2913 ( .IN1(g1027), .IN2(g1068), .S(n2007), .Q(g6894) );
  MUX21X1 U2914 ( .IN1(g1636), .IN2(n1969), .S(n2007), .Q(g8779) );
  AO21X1 U2915 ( .IN1(g554), .IN2(n1971), .IN3(n1970), .Q(g10793) );
  OA21X1 U2916 ( .IN1(n1973), .IN2(n1972), .IN3(n1997), .Q(n1974) );
  AO21X1 U2917 ( .IN1(n1998), .IN2(g1941), .IN3(n1974), .Q(n1975) );
  MUX21X1 U2918 ( .IN1(g1936), .IN2(n1976), .S(n1975), .Q(n1977) );
  AO21X1 U2919 ( .IN1(n2002), .IN2(n1977), .IN3(n1741), .Q(g8944) );
  MUX21X1 U2920 ( .IN1(n1979), .IN2(g1654), .S(n1978), .Q(g10765) );
  AO22X1 U2921 ( .IN1(g718), .IN2(n2004), .IN3(g727), .IN4(n2003), .Q(g8434)
         );
  MUX21X1 U2922 ( .IN1(g1453), .IN2(g1564), .S(n1992), .Q(g6546) );
  MUX21X1 U2923 ( .IN1(g148), .IN2(g269), .S(n2005), .Q(g6906) );
  INVX0 U2924 ( .INP(n1982), .ZN(g11324) );
  NAND2X0 U2925 ( .IN1(n1984), .IN2(n1983), .QN(n1987) );
  OA221X1 U2926 ( .IN1(n1987), .IN2(g673), .IN3(n1987), .IN4(n1986), .IN5(
        n1985), .Q(n1988) );
  MUX21X1 U2927 ( .IN1(g668), .IN2(n1807), .S(n1988), .Q(n1990) );
  AO21X1 U2928 ( .IN1(n1991), .IN2(n1990), .IN3(n1989), .Q(g8922) );
  MUX21X1 U2929 ( .IN1(g1515), .IN2(g1574), .S(n1992), .Q(g6478) );
  MUX21X1 U2930 ( .IN1(g131), .IN2(g290), .S(n2005), .Q(g6907) );
  INVX0 U2931 ( .INP(n1993), .ZN(n1994) );
  NAND2X0 U2932 ( .IN1(n1995), .IN2(n1994), .QN(n1996) );
  AO22X1 U2933 ( .IN1(n1998), .IN2(g1896), .IN3(n1997), .IN4(n1996), .Q(n1999)
         );
  MUX21X1 U2934 ( .IN1(g1891), .IN2(n2000), .S(n1999), .Q(n2001) );
  AO21X1 U2935 ( .IN1(n2002), .IN2(n2001), .IN3(n1741), .Q(g8937) );
  MUX21X1 U2936 ( .IN1(g158), .IN2(g275), .S(n2005), .Q(g6915) );
  AO22X1 U2937 ( .IN1(g700), .IN2(n2004), .IN3(g709), .IN4(n2003), .Q(g8432)
         );
  MUX21X1 U2938 ( .IN1(g174), .IN2(g281), .S(n2005), .Q(g6928) );
  MUX21X1 U2939 ( .IN1(g1015), .IN2(g1074), .S(n2007), .Q(g6930) );
  MUX21X1 U2940 ( .IN1(g1086), .IN2(g354), .S(n2006), .Q(g6071) );
  AO22X1 U2941 ( .IN1(n1289), .IN2(g1260), .IN3(g1265), .IN4(n1028), .Q(g7302)
         );
  MUX21X1 U2942 ( .IN1(g1007), .IN2(g1095), .S(n2007), .Q(g6918) );
  MUX21X1 U2943 ( .IN1(n1025), .IN2(g348), .S(n2008), .Q(g11481) );
  AO22X1 U2944 ( .IN1(n1289), .IN2(g1275), .IN3(g1235), .IN4(n1028), .Q(g7296)
         );
  XNOR2X1 U2945 ( .IN1(g590), .IN2(n2011), .Q(N599) );
  NOR2X0 U2946 ( .IN1(g1707), .IN2(n1008), .QN(g4076) );
  INVX0 U2947 ( .INP(g1707), .ZN(n2012) );
  OA221X1 U2948 ( .IN1(g1690), .IN2(g1707), .IN3(n2013), .IN4(n2012), .IN5(
        g1700), .Q(g6155) );
  OR3X1 U2949 ( .IN1(n2016), .IN2(n2015), .IN3(n2014), .Q(n2018) );
  NAND4X0 U2950 ( .IN1(g1690), .IN2(g1796), .IN3(g1806), .IN4(g1707), .QN(
        n2017) );
  NOR4X0 U2951 ( .IN1(g1781), .IN2(n2019), .IN3(n2018), .IN4(n2017), .QN(g5556) );
  AND2X1 U2952 ( .IN1(n2020), .IN2(g746), .Q(g2791) );
  AO22X1 U2953 ( .IN1(g754), .IN2(g2791), .IN3(n2021), .IN4(g746), .Q(g3462)
         );
  NAND2X0 U2954 ( .IN1(g109), .IN2(g108), .QN(n2022) );
  AND2X1 U2955 ( .IN1(n2023), .IN2(n2022), .Q(g5763) );
  INVX0 U2956 ( .INP(g23), .ZN(g3327) );
  INVX0 U2957 ( .INP(n2024), .ZN(n2025) );
  NOR2X0 U2958 ( .IN1(g32), .IN2(n2025), .QN(n2027) );
  XNOR2X1 U2959 ( .IN1(n2027), .IN2(n2026), .Q(g11286) );
  XOR2X1 U2960 ( .IN1(n2028), .IN2(g11286), .Q(g11163) );
endmodule

